module AXI4StreamToBundleBridge(
  output        auto_in_ready,
  input         auto_in_valid,
  input  [63:0] auto_in_bits_data,
  input         auto_in_bits_last,
  input         auto_out_ready,
  output        auto_out_valid,
  output [63:0] auto_out_bits_data,
  output        auto_out_bits_last
);
  assign auto_in_ready = auto_out_ready; // @[LazyModule.scala 173:31]
  assign auto_out_valid = auto_in_valid; // @[LazyModule.scala 173:49]
  assign auto_out_bits_data = auto_in_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_bits_last = auto_in_bits_last; // @[LazyModule.scala 173:49]
endmodule
module ConstantCoefficientFIRFilter(
  input         clock,
  input         reset,
  input         io_in_valid,
  input  [31:0] io_in_bits,
  output        io_out_valid,
  output [31:0] io_out_bits
);
  reg [31:0] regs_0; // @[FIRFilter.scala 39:21]
  reg [31:0] _RAND_0;
  reg [31:0] regs_1; // @[FIRFilter.scala 39:21]
  reg [31:0] _RAND_1;
  reg [31:0] regs_2; // @[FIRFilter.scala 39:21]
  reg [31:0] _RAND_2;
  reg [31:0] regs_3; // @[FIRFilter.scala 39:21]
  reg [31:0] _RAND_3;
  reg [31:0] regs_4; // @[FIRFilter.scala 39:21]
  reg [31:0] _RAND_4;
  reg [31:0] regs_5; // @[FIRFilter.scala 39:21]
  reg [31:0] _RAND_5;
  wire [47:0] accumulator_0; // @[FixedPointTypeClass.scala 43:59]
  wire [48:0] muls_1; // @[FixedPointTypeClass.scala 43:59]
  wire [48:0] muls_2; // @[FixedPointTypeClass.scala 43:59]
  wire [49:0] muls_3; // @[FixedPointTypeClass.scala 43:59]
  wire [49:0] muls_4; // @[FixedPointTypeClass.scala 43:59]
  wire [32:0] muls_5; // @[FixedPointTypeClass.scala 43:59]
  wire [48:0] _GEN_19; // @[FixedPointTypeClass.scala 21:58]
  wire [48:0] _T_8; // @[FixedPointTypeClass.scala 21:58]
  wire [48:0] accumulator_1; // @[FixedPointTypeClass.scala 21:58]
  wire [48:0] _T_10; // @[FixedPointTypeClass.scala 21:58]
  wire [48:0] accumulator_2; // @[FixedPointTypeClass.scala 21:58]
  wire [49:0] _GEN_20; // @[FixedPointTypeClass.scala 21:58]
  wire [49:0] _T_12; // @[FixedPointTypeClass.scala 21:58]
  wire [49:0] accumulator_3; // @[FixedPointTypeClass.scala 21:58]
  wire [49:0] _T_14; // @[FixedPointTypeClass.scala 21:58]
  wire [49:0] accumulator_4; // @[FixedPointTypeClass.scala 21:58]
  wire [49:0] _GEN_21; // @[FixedPointTypeClass.scala 21:58]
  wire [49:0] _T_16; // @[FixedPointTypeClass.scala 21:58]
  wire [49:0] accumulator_5; // @[FixedPointTypeClass.scala 21:58]
  reg  _T_18; // @[Reg.scala 19:20]
  reg [31:0] _RAND_6;
  reg  _T_19; // @[Reg.scala 19:20]
  reg [31:0] _RAND_7;
  reg  _T_20; // @[Reg.scala 19:20]
  reg [31:0] _RAND_8;
  reg  _T_21; // @[Reg.scala 19:20]
  reg [31:0] _RAND_9;
  reg  _T_22; // @[Reg.scala 19:20]
  reg [31:0] _RAND_10;
  reg  _T_23; // @[Reg.scala 19:20]
  reg [31:0] _RAND_11;
  wire [35:0] _GEN_22; // @[FIRFilter.scala 67:15]
  wire [31:0] _GEN_23; // @[FIRFilter.scala 67:15]
  assign accumulator_0 = $signed(regs_0) * $signed(32'sh4000); // @[FixedPointTypeClass.scala 43:59]
  assign muls_1 = $signed(regs_1) * $signed(32'sh8000); // @[FixedPointTypeClass.scala 43:59]
  assign muls_2 = $signed(regs_2) * $signed(32'shc000); // @[FixedPointTypeClass.scala 43:59]
  assign muls_3 = $signed(regs_3) * $signed(32'sh10000); // @[FixedPointTypeClass.scala 43:59]
  assign muls_4 = $signed(regs_4) * $signed(32'sh14000); // @[FixedPointTypeClass.scala 43:59]
  assign muls_5 = $signed(regs_5) * $signed(32'sh0); // @[FixedPointTypeClass.scala 43:59]
  assign _GEN_19 = {{1{accumulator_0[47]}},accumulator_0}; // @[FixedPointTypeClass.scala 21:58]
  assign _T_8 = $signed(muls_1) + $signed(_GEN_19); // @[FixedPointTypeClass.scala 21:58]
  assign accumulator_1 = $signed(_T_8); // @[FixedPointTypeClass.scala 21:58]
  assign _T_10 = $signed(muls_2) + $signed(accumulator_1); // @[FixedPointTypeClass.scala 21:58]
  assign accumulator_2 = $signed(_T_10); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_20 = {{1{accumulator_2[48]}},accumulator_2}; // @[FixedPointTypeClass.scala 21:58]
  assign _T_12 = $signed(muls_3) + $signed(_GEN_20); // @[FixedPointTypeClass.scala 21:58]
  assign accumulator_3 = $signed(_T_12); // @[FixedPointTypeClass.scala 21:58]
  assign _T_14 = $signed(muls_4) + $signed(accumulator_3); // @[FixedPointTypeClass.scala 21:58]
  assign accumulator_4 = $signed(_T_14); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_21 = {{17{muls_5[32]}},muls_5}; // @[FixedPointTypeClass.scala 21:58]
  assign _T_16 = $signed(_GEN_21) + $signed(accumulator_4); // @[FixedPointTypeClass.scala 21:58]
  assign accumulator_5 = $signed(_T_16); // @[FixedPointTypeClass.scala 21:58]
  assign io_out_valid = _T_23 & io_in_valid; // @[FIRFilter.scala 68:16]
  assign _GEN_22 = accumulator_5[49:14]; // @[FIRFilter.scala 67:15]
  assign _GEN_23 = _GEN_22[31:0]; // @[FIRFilter.scala 67:15]
  assign io_out_bits = $signed(_GEN_23); // @[FIRFilter.scala 67:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  regs_3 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  regs_4 = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  regs_5 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_18 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_19 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_20 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_21 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_22 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_23 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      regs_0 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_0 <= io_in_bits;
      end
    end
    if (reset) begin
      regs_1 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_1 <= regs_0;
      end
    end
    if (reset) begin
      regs_2 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_2 <= regs_1;
      end
    end
    if (reset) begin
      regs_3 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_3 <= regs_2;
      end
    end
    if (reset) begin
      regs_4 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_4 <= regs_3;
      end
    end
    if (reset) begin
      regs_5 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_5 <= regs_4;
      end
    end
    if (reset) begin
      _T_18 <= 1'h0;
    end else begin
      if (io_in_valid) begin
        _T_18 <= io_in_valid;
      end
    end
    if (reset) begin
      _T_19 <= 1'h0;
    end else begin
      if (io_in_valid) begin
        _T_19 <= _T_18;
      end
    end
    if (reset) begin
      _T_20 <= 1'h0;
    end else begin
      if (io_in_valid) begin
        _T_20 <= _T_19;
      end
    end
    if (reset) begin
      _T_21 <= 1'h0;
    end else begin
      if (io_in_valid) begin
        _T_21 <= _T_20;
      end
    end
    if (reset) begin
      _T_22 <= 1'h0;
    end else begin
      if (io_in_valid) begin
        _T_22 <= _T_21;
      end
    end
    if (reset) begin
      _T_23 <= 1'h0;
    end else begin
      if (io_in_valid) begin
        _T_23 <= _T_22;
      end
    end
  end
endmodule
module lineLength(
  input         clock,
  input         reset,
  input         io_in_valid,
  input  [31:0] io_in_bits,
  output        io_out_valid,
  output [31:0] io_out_bits
);
  reg [31:0] lineLengths_0; // @[lineLength.scala 47:28]
  reg [31:0] _RAND_0;
  reg [31:0] pastVal; // @[lineLength.scala 49:24]
  reg [31:0] _RAND_1;
  wire  _T_3; // @[FixedPointTypeClass.scala 57:62]
  wire [31:0] _T_5; // @[FixedPointTypeClass.scala 31:68]
  wire [31:0] _T_6; // @[FixedPointTypeClass.scala 31:68]
  wire [31:0] _T_8; // @[FixedPointTypeClass.scala 31:68]
  wire [31:0] _T_9; // @[FixedPointTypeClass.scala 31:68]
  wire [30:0] _T_12; // @[FixedPointTypeClass.scala 118:50]
  wire [27:0] _T_13; // @[FixedPointTypeClass.scala 118:50]
  reg  _T_14; // @[Reg.scala 19:20]
  reg [31:0] _RAND_2;
  reg  _T_15; // @[Reg.scala 19:20]
  reg [31:0] _RAND_3;
  assign _T_3 = $signed(io_in_bits) >= $signed(pastVal); // @[FixedPointTypeClass.scala 57:62]
  assign _T_5 = $signed(io_in_bits) - $signed(pastVal); // @[FixedPointTypeClass.scala 31:68]
  assign _T_6 = $signed(_T_5); // @[FixedPointTypeClass.scala 31:68]
  assign _T_8 = $signed(pastVal) - $signed(io_in_bits); // @[FixedPointTypeClass.scala 31:68]
  assign _T_9 = $signed(_T_8); // @[FixedPointTypeClass.scala 31:68]
  assign _T_12 = lineLengths_0[31:1]; // @[FixedPointTypeClass.scala 118:50]
  assign _T_13 = _T_12[30:3]; // @[FixedPointTypeClass.scala 118:50]
  assign io_out_valid = _T_15 & io_in_valid; // @[lineLength.scala 84:16]
  assign io_out_bits = {{4{_T_13[27]}},_T_13}; // @[lineLength.scala 83:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  lineLengths_0 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  pastVal = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_14 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_15 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      lineLengths_0 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        if (_T_3) begin
          lineLengths_0 <= _T_6;
        end else begin
          lineLengths_0 <= _T_9;
        end
      end
    end
    if (reset) begin
      pastVal <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        pastVal <= io_in_bits;
      end
    end
    if (reset) begin
      _T_14 <= 1'h0;
    end else begin
      if (io_in_valid) begin
        _T_14 <= io_in_valid;
      end
    end
    if (reset) begin
      _T_15 <= 1'h0;
    end else begin
      if (io_in_valid) begin
        _T_15 <= _T_14;
      end
    end
  end
endmodule
module sumSquares(
  input         clock,
  input         reset,
  input         io_in_valid,
  input  [31:0] io_in_bits,
  output        io_out_valid,
  output [31:0] io_out_bits
);
  reg [31:0] sumSquaress_0; // @[SumSquares.scala 41:28]
  reg [31:0] _RAND_0;
  wire [63:0] _T_3; // @[FixedPointTypeClass.scala 43:59]
  wire [39:0] _GEN_7; // @[SumSquares.scala 52:31]
  wire [39:0] _GEN_8; // @[SumSquares.scala 52:31]
  wire [63:0] _GEN_1; // @[SumSquares.scala 52:31]
  wire [30:0] _T_5; // @[FixedPointTypeClass.scala 118:50]
  wire [27:0] _T_6; // @[FixedPointTypeClass.scala 118:50]
  reg  _T_7; // @[Reg.scala 19:20]
  reg [31:0] _RAND_1;
  reg  _T_8; // @[Reg.scala 19:20]
  reg [31:0] _RAND_2;
  wire [55:0] _GEN_10; // @[SumSquares.scala 53:34 SumSquares.scala 56:22]
  wire [31:0] _GEN_11; // @[SumSquares.scala 53:34 SumSquares.scala 56:22]
  assign _T_3 = $signed(io_in_bits) * $signed(io_in_bits); // @[FixedPointTypeClass.scala 43:59]
  assign _GEN_7 = {{8{sumSquaress_0[31]}},sumSquaress_0}; // @[SumSquares.scala 52:31]
  assign _GEN_8 = $signed(_GEN_7) << 8; // @[SumSquares.scala 52:31]
  assign _GEN_1 = io_in_valid ? $signed(_T_3) : $signed({{24{_GEN_8[39]}},_GEN_8}); // @[SumSquares.scala 52:31]
  assign _T_5 = sumSquaress_0[31:1]; // @[FixedPointTypeClass.scala 118:50]
  assign _T_6 = _T_5[30:3]; // @[FixedPointTypeClass.scala 118:50]
  assign io_out_valid = _T_8 & io_in_valid; // @[SumSquares.scala 78:16]
  assign io_out_bits = {{4{_T_6[27]}},_T_6}; // @[SumSquares.scala 77:15]
  assign _GEN_10 = _GEN_1[63:8]; // @[SumSquares.scala 53:34 SumSquares.scala 56:22]
  assign _GEN_11 = _GEN_10[31:0]; // @[SumSquares.scala 53:34 SumSquares.scala 56:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sumSquaress_0 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_7 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_8 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      sumSquaress_0 <= 32'sh0;
    end else begin
      sumSquaress_0 <= $signed(_GEN_11);
    end
    if (reset) begin
      _T_7 <= 1'h0;
    end else begin
      if (io_in_valid) begin
        _T_7 <= io_in_valid;
      end
    end
    if (reset) begin
      _T_8 <= 1'h0;
    end else begin
      if (io_in_valid) begin
        _T_8 <= _T_7;
      end
    end
  end
endmodule
module NeuralNet(
  input         clock,
  input         io_in_valid,
  input  [31:0] io_in_bits_0,
  input  [31:0] io_in_bits_1,
  input  [31:0] io_in_bits_2,
  input  [31:0] io_in_bits_3,
  output        io_out_valid,
  output        io_out_bits,
  input  [31:0] io_weightMatrix_0_0,
  input  [31:0] io_weightMatrix_0_1,
  input  [31:0] io_weightMatrix_0_2,
  input  [31:0] io_weightMatrix_0_3,
  input  [31:0] io_weightMatrix_1_0,
  input  [31:0] io_weightMatrix_1_1,
  input  [31:0] io_weightMatrix_1_2,
  input  [31:0] io_weightMatrix_1_3,
  input  [31:0] io_weightMatrix_2_0,
  input  [31:0] io_weightMatrix_2_1,
  input  [31:0] io_weightMatrix_2_2,
  input  [31:0] io_weightMatrix_2_3,
  input  [31:0] io_weightMatrix_3_0,
  input  [31:0] io_weightMatrix_3_1,
  input  [31:0] io_weightMatrix_3_2,
  input  [31:0] io_weightMatrix_3_3,
  input  [31:0] io_weightMatrix_4_0,
  input  [31:0] io_weightMatrix_4_1,
  input  [31:0] io_weightMatrix_4_2,
  input  [31:0] io_weightMatrix_4_3,
  input  [31:0] io_weightMatrix_5_0,
  input  [31:0] io_weightMatrix_5_1,
  input  [31:0] io_weightMatrix_5_2,
  input  [31:0] io_weightMatrix_5_3,
  input  [31:0] io_weightMatrix_6_0,
  input  [31:0] io_weightMatrix_6_1,
  input  [31:0] io_weightMatrix_6_2,
  input  [31:0] io_weightMatrix_6_3,
  input  [31:0] io_weightMatrix_7_0,
  input  [31:0] io_weightMatrix_7_1,
  input  [31:0] io_weightMatrix_7_2,
  input  [31:0] io_weightMatrix_7_3,
  input  [31:0] io_weightMatrix_8_0,
  input  [31:0] io_weightMatrix_8_1,
  input  [31:0] io_weightMatrix_8_2,
  input  [31:0] io_weightMatrix_8_3,
  input  [31:0] io_weightMatrix_9_0,
  input  [31:0] io_weightMatrix_9_1,
  input  [31:0] io_weightMatrix_9_2,
  input  [31:0] io_weightMatrix_9_3,
  input  [31:0] io_weightMatrix_10_0,
  input  [31:0] io_weightMatrix_10_1,
  input  [31:0] io_weightMatrix_10_2,
  input  [31:0] io_weightMatrix_10_3,
  input  [31:0] io_weightMatrix_11_0,
  input  [31:0] io_weightMatrix_11_1,
  input  [31:0] io_weightMatrix_11_2,
  input  [31:0] io_weightMatrix_11_3,
  input  [31:0] io_weightMatrix_12_0,
  input  [31:0] io_weightMatrix_12_1,
  input  [31:0] io_weightMatrix_12_2,
  input  [31:0] io_weightMatrix_12_3,
  input  [31:0] io_weightMatrix_13_0,
  input  [31:0] io_weightMatrix_13_1,
  input  [31:0] io_weightMatrix_13_2,
  input  [31:0] io_weightMatrix_13_3,
  input  [31:0] io_weightMatrix_14_0,
  input  [31:0] io_weightMatrix_14_1,
  input  [31:0] io_weightMatrix_14_2,
  input  [31:0] io_weightMatrix_14_3,
  input  [31:0] io_weightMatrix_15_0,
  input  [31:0] io_weightMatrix_15_1,
  input  [31:0] io_weightMatrix_15_2,
  input  [31:0] io_weightMatrix_15_3,
  input  [31:0] io_weightMatrix_16_0,
  input  [31:0] io_weightMatrix_16_1,
  input  [31:0] io_weightMatrix_16_2,
  input  [31:0] io_weightMatrix_16_3,
  input  [31:0] io_weightMatrix_17_0,
  input  [31:0] io_weightMatrix_17_1,
  input  [31:0] io_weightMatrix_17_2,
  input  [31:0] io_weightMatrix_17_3,
  input  [31:0] io_weightMatrix_18_0,
  input  [31:0] io_weightMatrix_18_1,
  input  [31:0] io_weightMatrix_18_2,
  input  [31:0] io_weightMatrix_18_3,
  input  [31:0] io_weightMatrix_19_0,
  input  [31:0] io_weightMatrix_19_1,
  input  [31:0] io_weightMatrix_19_2,
  input  [31:0] io_weightMatrix_19_3,
  input  [31:0] io_weightMatrix_20_0,
  input  [31:0] io_weightMatrix_20_1,
  input  [31:0] io_weightMatrix_20_2,
  input  [31:0] io_weightMatrix_20_3,
  input  [31:0] io_weightMatrix_21_0,
  input  [31:0] io_weightMatrix_21_1,
  input  [31:0] io_weightMatrix_21_2,
  input  [31:0] io_weightMatrix_21_3,
  input  [31:0] io_weightMatrix_22_0,
  input  [31:0] io_weightMatrix_22_1,
  input  [31:0] io_weightMatrix_22_2,
  input  [31:0] io_weightMatrix_22_3,
  input  [31:0] io_weightMatrix_23_0,
  input  [31:0] io_weightMatrix_23_1,
  input  [31:0] io_weightMatrix_23_2,
  input  [31:0] io_weightMatrix_23_3,
  input  [31:0] io_weightMatrix_24_0,
  input  [31:0] io_weightMatrix_24_1,
  input  [31:0] io_weightMatrix_24_2,
  input  [31:0] io_weightMatrix_24_3,
  input  [31:0] io_weightMatrix_25_0,
  input  [31:0] io_weightMatrix_25_1,
  input  [31:0] io_weightMatrix_25_2,
  input  [31:0] io_weightMatrix_25_3,
  input  [31:0] io_weightMatrix_26_0,
  input  [31:0] io_weightMatrix_26_1,
  input  [31:0] io_weightMatrix_26_2,
  input  [31:0] io_weightMatrix_26_3,
  input  [31:0] io_weightMatrix_27_0,
  input  [31:0] io_weightMatrix_27_1,
  input  [31:0] io_weightMatrix_27_2,
  input  [31:0] io_weightMatrix_27_3,
  input  [31:0] io_weightMatrix_28_0,
  input  [31:0] io_weightMatrix_28_1,
  input  [31:0] io_weightMatrix_28_2,
  input  [31:0] io_weightMatrix_28_3,
  input  [31:0] io_weightMatrix_29_0,
  input  [31:0] io_weightMatrix_29_1,
  input  [31:0] io_weightMatrix_29_2,
  input  [31:0] io_weightMatrix_29_3,
  input  [31:0] io_weightMatrix_30_0,
  input  [31:0] io_weightMatrix_30_1,
  input  [31:0] io_weightMatrix_30_2,
  input  [31:0] io_weightMatrix_30_3,
  input  [31:0] io_weightMatrix_31_0,
  input  [31:0] io_weightMatrix_31_1,
  input  [31:0] io_weightMatrix_31_2,
  input  [31:0] io_weightMatrix_31_3,
  input  [31:0] io_weightMatrix_32_0,
  input  [31:0] io_weightMatrix_32_1,
  input  [31:0] io_weightMatrix_32_2,
  input  [31:0] io_weightMatrix_32_3,
  input  [31:0] io_weightMatrix_33_0,
  input  [31:0] io_weightMatrix_33_1,
  input  [31:0] io_weightMatrix_33_2,
  input  [31:0] io_weightMatrix_33_3,
  input  [31:0] io_weightMatrix_34_0,
  input  [31:0] io_weightMatrix_34_1,
  input  [31:0] io_weightMatrix_34_2,
  input  [31:0] io_weightMatrix_34_3,
  input  [31:0] io_weightMatrix_35_0,
  input  [31:0] io_weightMatrix_35_1,
  input  [31:0] io_weightMatrix_35_2,
  input  [31:0] io_weightMatrix_35_3,
  input  [31:0] io_weightMatrix_36_0,
  input  [31:0] io_weightMatrix_36_1,
  input  [31:0] io_weightMatrix_36_2,
  input  [31:0] io_weightMatrix_36_3,
  input  [31:0] io_weightMatrix_37_0,
  input  [31:0] io_weightMatrix_37_1,
  input  [31:0] io_weightMatrix_37_2,
  input  [31:0] io_weightMatrix_37_3,
  input  [31:0] io_weightMatrix_38_0,
  input  [31:0] io_weightMatrix_38_1,
  input  [31:0] io_weightMatrix_38_2,
  input  [31:0] io_weightMatrix_38_3,
  input  [31:0] io_weightMatrix_39_0,
  input  [31:0] io_weightMatrix_39_1,
  input  [31:0] io_weightMatrix_39_2,
  input  [31:0] io_weightMatrix_39_3,
  input  [31:0] io_weightMatrix_40_0,
  input  [31:0] io_weightMatrix_40_1,
  input  [31:0] io_weightMatrix_40_2,
  input  [31:0] io_weightMatrix_40_3,
  input  [31:0] io_weightMatrix_41_0,
  input  [31:0] io_weightMatrix_41_1,
  input  [31:0] io_weightMatrix_41_2,
  input  [31:0] io_weightMatrix_41_3,
  input  [31:0] io_weightMatrix_42_0,
  input  [31:0] io_weightMatrix_42_1,
  input  [31:0] io_weightMatrix_42_2,
  input  [31:0] io_weightMatrix_42_3,
  input  [31:0] io_weightMatrix_43_0,
  input  [31:0] io_weightMatrix_43_1,
  input  [31:0] io_weightMatrix_43_2,
  input  [31:0] io_weightMatrix_43_3,
  input  [31:0] io_weightMatrix_44_0,
  input  [31:0] io_weightMatrix_44_1,
  input  [31:0] io_weightMatrix_44_2,
  input  [31:0] io_weightMatrix_44_3,
  input  [31:0] io_weightMatrix_45_0,
  input  [31:0] io_weightMatrix_45_1,
  input  [31:0] io_weightMatrix_45_2,
  input  [31:0] io_weightMatrix_45_3,
  input  [31:0] io_weightMatrix_46_0,
  input  [31:0] io_weightMatrix_46_1,
  input  [31:0] io_weightMatrix_46_2,
  input  [31:0] io_weightMatrix_46_3,
  input  [31:0] io_weightMatrix_47_0,
  input  [31:0] io_weightMatrix_47_1,
  input  [31:0] io_weightMatrix_47_2,
  input  [31:0] io_weightMatrix_47_3,
  input  [31:0] io_weightMatrix_48_0,
  input  [31:0] io_weightMatrix_48_1,
  input  [31:0] io_weightMatrix_48_2,
  input  [31:0] io_weightMatrix_48_3,
  input  [31:0] io_weightMatrix_49_0,
  input  [31:0] io_weightMatrix_49_1,
  input  [31:0] io_weightMatrix_49_2,
  input  [31:0] io_weightMatrix_49_3,
  input  [31:0] io_weightMatrix_50_0,
  input  [31:0] io_weightMatrix_50_1,
  input  [31:0] io_weightMatrix_50_2,
  input  [31:0] io_weightMatrix_50_3,
  input  [31:0] io_weightMatrix_51_0,
  input  [31:0] io_weightMatrix_51_1,
  input  [31:0] io_weightMatrix_51_2,
  input  [31:0] io_weightMatrix_51_3,
  input  [31:0] io_weightMatrix_52_0,
  input  [31:0] io_weightMatrix_52_1,
  input  [31:0] io_weightMatrix_52_2,
  input  [31:0] io_weightMatrix_52_3,
  input  [31:0] io_weightMatrix_53_0,
  input  [31:0] io_weightMatrix_53_1,
  input  [31:0] io_weightMatrix_53_2,
  input  [31:0] io_weightMatrix_53_3,
  input  [31:0] io_weightMatrix_54_0,
  input  [31:0] io_weightMatrix_54_1,
  input  [31:0] io_weightMatrix_54_2,
  input  [31:0] io_weightMatrix_54_3,
  input  [31:0] io_weightMatrix_55_0,
  input  [31:0] io_weightMatrix_55_1,
  input  [31:0] io_weightMatrix_55_2,
  input  [31:0] io_weightMatrix_55_3,
  input  [31:0] io_weightMatrix_56_0,
  input  [31:0] io_weightMatrix_56_1,
  input  [31:0] io_weightMatrix_56_2,
  input  [31:0] io_weightMatrix_56_3,
  input  [31:0] io_weightMatrix_57_0,
  input  [31:0] io_weightMatrix_57_1,
  input  [31:0] io_weightMatrix_57_2,
  input  [31:0] io_weightMatrix_57_3,
  input  [31:0] io_weightMatrix_58_0,
  input  [31:0] io_weightMatrix_58_1,
  input  [31:0] io_weightMatrix_58_2,
  input  [31:0] io_weightMatrix_58_3,
  input  [31:0] io_weightMatrix_59_0,
  input  [31:0] io_weightMatrix_59_1,
  input  [31:0] io_weightMatrix_59_2,
  input  [31:0] io_weightMatrix_59_3,
  input  [31:0] io_weightMatrix_60_0,
  input  [31:0] io_weightMatrix_60_1,
  input  [31:0] io_weightMatrix_60_2,
  input  [31:0] io_weightMatrix_60_3,
  input  [31:0] io_weightMatrix_61_0,
  input  [31:0] io_weightMatrix_61_1,
  input  [31:0] io_weightMatrix_61_2,
  input  [31:0] io_weightMatrix_61_3,
  input  [31:0] io_weightMatrix_62_0,
  input  [31:0] io_weightMatrix_62_1,
  input  [31:0] io_weightMatrix_62_2,
  input  [31:0] io_weightMatrix_62_3,
  input  [31:0] io_weightMatrix_63_0,
  input  [31:0] io_weightMatrix_63_1,
  input  [31:0] io_weightMatrix_63_2,
  input  [31:0] io_weightMatrix_63_3,
  input  [31:0] io_weightMatrix_64_0,
  input  [31:0] io_weightMatrix_64_1,
  input  [31:0] io_weightMatrix_64_2,
  input  [31:0] io_weightMatrix_64_3,
  input  [31:0] io_weightMatrix_65_0,
  input  [31:0] io_weightMatrix_65_1,
  input  [31:0] io_weightMatrix_65_2,
  input  [31:0] io_weightMatrix_65_3,
  input  [31:0] io_weightMatrix_66_0,
  input  [31:0] io_weightMatrix_66_1,
  input  [31:0] io_weightMatrix_66_2,
  input  [31:0] io_weightMatrix_66_3,
  input  [31:0] io_weightMatrix_67_0,
  input  [31:0] io_weightMatrix_67_1,
  input  [31:0] io_weightMatrix_67_2,
  input  [31:0] io_weightMatrix_67_3,
  input  [31:0] io_weightMatrix_68_0,
  input  [31:0] io_weightMatrix_68_1,
  input  [31:0] io_weightMatrix_68_2,
  input  [31:0] io_weightMatrix_68_3,
  input  [31:0] io_weightMatrix_69_0,
  input  [31:0] io_weightMatrix_69_1,
  input  [31:0] io_weightMatrix_69_2,
  input  [31:0] io_weightMatrix_69_3,
  input  [31:0] io_weightMatrix_70_0,
  input  [31:0] io_weightMatrix_70_1,
  input  [31:0] io_weightMatrix_70_2,
  input  [31:0] io_weightMatrix_70_3,
  input  [31:0] io_weightMatrix_71_0,
  input  [31:0] io_weightMatrix_71_1,
  input  [31:0] io_weightMatrix_71_2,
  input  [31:0] io_weightMatrix_71_3,
  input  [31:0] io_weightMatrix_72_0,
  input  [31:0] io_weightMatrix_72_1,
  input  [31:0] io_weightMatrix_72_2,
  input  [31:0] io_weightMatrix_72_3,
  input  [31:0] io_weightMatrix_73_0,
  input  [31:0] io_weightMatrix_73_1,
  input  [31:0] io_weightMatrix_73_2,
  input  [31:0] io_weightMatrix_73_3,
  input  [31:0] io_weightMatrix_74_0,
  input  [31:0] io_weightMatrix_74_1,
  input  [31:0] io_weightMatrix_74_2,
  input  [31:0] io_weightMatrix_74_3,
  input  [31:0] io_weightMatrix_75_0,
  input  [31:0] io_weightMatrix_75_1,
  input  [31:0] io_weightMatrix_75_2,
  input  [31:0] io_weightMatrix_75_3,
  input  [31:0] io_weightMatrix_76_0,
  input  [31:0] io_weightMatrix_76_1,
  input  [31:0] io_weightMatrix_76_2,
  input  [31:0] io_weightMatrix_76_3,
  input  [31:0] io_weightMatrix_77_0,
  input  [31:0] io_weightMatrix_77_1,
  input  [31:0] io_weightMatrix_77_2,
  input  [31:0] io_weightMatrix_77_3,
  input  [31:0] io_weightMatrix_78_0,
  input  [31:0] io_weightMatrix_78_1,
  input  [31:0] io_weightMatrix_78_2,
  input  [31:0] io_weightMatrix_78_3,
  input  [31:0] io_weightMatrix_79_0,
  input  [31:0] io_weightMatrix_79_1,
  input  [31:0] io_weightMatrix_79_2,
  input  [31:0] io_weightMatrix_79_3,
  input  [31:0] io_weightMatrix_80_0,
  input  [31:0] io_weightMatrix_80_1,
  input  [31:0] io_weightMatrix_80_2,
  input  [31:0] io_weightMatrix_80_3,
  input  [31:0] io_weightMatrix_81_0,
  input  [31:0] io_weightMatrix_81_1,
  input  [31:0] io_weightMatrix_81_2,
  input  [31:0] io_weightMatrix_81_3,
  input  [31:0] io_weightMatrix_82_0,
  input  [31:0] io_weightMatrix_82_1,
  input  [31:0] io_weightMatrix_82_2,
  input  [31:0] io_weightMatrix_82_3,
  input  [31:0] io_weightMatrix_83_0,
  input  [31:0] io_weightMatrix_83_1,
  input  [31:0] io_weightMatrix_83_2,
  input  [31:0] io_weightMatrix_83_3,
  input  [31:0] io_weightMatrix_84_0,
  input  [31:0] io_weightMatrix_84_1,
  input  [31:0] io_weightMatrix_84_2,
  input  [31:0] io_weightMatrix_84_3,
  input  [31:0] io_weightMatrix_85_0,
  input  [31:0] io_weightMatrix_85_1,
  input  [31:0] io_weightMatrix_85_2,
  input  [31:0] io_weightMatrix_85_3,
  input  [31:0] io_weightMatrix_86_0,
  input  [31:0] io_weightMatrix_86_1,
  input  [31:0] io_weightMatrix_86_2,
  input  [31:0] io_weightMatrix_86_3,
  input  [31:0] io_weightMatrix_87_0,
  input  [31:0] io_weightMatrix_87_1,
  input  [31:0] io_weightMatrix_87_2,
  input  [31:0] io_weightMatrix_87_3,
  input  [31:0] io_weightMatrix_88_0,
  input  [31:0] io_weightMatrix_88_1,
  input  [31:0] io_weightMatrix_88_2,
  input  [31:0] io_weightMatrix_88_3,
  input  [31:0] io_weightMatrix_89_0,
  input  [31:0] io_weightMatrix_89_1,
  input  [31:0] io_weightMatrix_89_2,
  input  [31:0] io_weightMatrix_89_3,
  input  [31:0] io_weightMatrix_90_0,
  input  [31:0] io_weightMatrix_90_1,
  input  [31:0] io_weightMatrix_90_2,
  input  [31:0] io_weightMatrix_90_3,
  input  [31:0] io_weightMatrix_91_0,
  input  [31:0] io_weightMatrix_91_1,
  input  [31:0] io_weightMatrix_91_2,
  input  [31:0] io_weightMatrix_91_3,
  input  [31:0] io_weightMatrix_92_0,
  input  [31:0] io_weightMatrix_92_1,
  input  [31:0] io_weightMatrix_92_2,
  input  [31:0] io_weightMatrix_92_3,
  input  [31:0] io_weightMatrix_93_0,
  input  [31:0] io_weightMatrix_93_1,
  input  [31:0] io_weightMatrix_93_2,
  input  [31:0] io_weightMatrix_93_3,
  input  [31:0] io_weightMatrix_94_0,
  input  [31:0] io_weightMatrix_94_1,
  input  [31:0] io_weightMatrix_94_2,
  input  [31:0] io_weightMatrix_94_3,
  input  [31:0] io_weightMatrix_95_0,
  input  [31:0] io_weightMatrix_95_1,
  input  [31:0] io_weightMatrix_95_2,
  input  [31:0] io_weightMatrix_95_3,
  input  [31:0] io_weightMatrix_96_0,
  input  [31:0] io_weightMatrix_96_1,
  input  [31:0] io_weightMatrix_96_2,
  input  [31:0] io_weightMatrix_96_3,
  input  [31:0] io_weightMatrix_97_0,
  input  [31:0] io_weightMatrix_97_1,
  input  [31:0] io_weightMatrix_97_2,
  input  [31:0] io_weightMatrix_97_3,
  input  [31:0] io_weightMatrix_98_0,
  input  [31:0] io_weightMatrix_98_1,
  input  [31:0] io_weightMatrix_98_2,
  input  [31:0] io_weightMatrix_98_3,
  input  [31:0] io_weightMatrix_99_0,
  input  [31:0] io_weightMatrix_99_1,
  input  [31:0] io_weightMatrix_99_2,
  input  [31:0] io_weightMatrix_99_3,
  input  [31:0] io_weightVec_0,
  input  [31:0] io_weightVec_1,
  input  [31:0] io_weightVec_2,
  input  [31:0] io_weightVec_3,
  input  [31:0] io_weightVec_4,
  input  [31:0] io_weightVec_5,
  input  [31:0] io_weightVec_6,
  input  [31:0] io_weightVec_7,
  input  [31:0] io_weightVec_8,
  input  [31:0] io_weightVec_9,
  input  [31:0] io_weightVec_10,
  input  [31:0] io_weightVec_11,
  input  [31:0] io_weightVec_12,
  input  [31:0] io_weightVec_13,
  input  [31:0] io_weightVec_14,
  input  [31:0] io_weightVec_15,
  input  [31:0] io_weightVec_16,
  input  [31:0] io_weightVec_17,
  input  [31:0] io_weightVec_18,
  input  [31:0] io_weightVec_19,
  input  [31:0] io_weightVec_20,
  input  [31:0] io_weightVec_21,
  input  [31:0] io_weightVec_22,
  input  [31:0] io_weightVec_23,
  input  [31:0] io_weightVec_24,
  input  [31:0] io_weightVec_25,
  input  [31:0] io_weightVec_26,
  input  [31:0] io_weightVec_27,
  input  [31:0] io_weightVec_28,
  input  [31:0] io_weightVec_29,
  input  [31:0] io_weightVec_30,
  input  [31:0] io_weightVec_31,
  input  [31:0] io_weightVec_32,
  input  [31:0] io_weightVec_33,
  input  [31:0] io_weightVec_34,
  input  [31:0] io_weightVec_35,
  input  [31:0] io_weightVec_36,
  input  [31:0] io_weightVec_37,
  input  [31:0] io_weightVec_38,
  input  [31:0] io_weightVec_39,
  input  [31:0] io_weightVec_40,
  input  [31:0] io_weightVec_41,
  input  [31:0] io_weightVec_42,
  input  [31:0] io_weightVec_43,
  input  [31:0] io_weightVec_44,
  input  [31:0] io_weightVec_45,
  input  [31:0] io_weightVec_46,
  input  [31:0] io_weightVec_47,
  input  [31:0] io_weightVec_48,
  input  [31:0] io_weightVec_49,
  input  [31:0] io_weightVec_50,
  input  [31:0] io_weightVec_51,
  input  [31:0] io_weightVec_52,
  input  [31:0] io_weightVec_53,
  input  [31:0] io_weightVec_54,
  input  [31:0] io_weightVec_55,
  input  [31:0] io_weightVec_56,
  input  [31:0] io_weightVec_57,
  input  [31:0] io_weightVec_58,
  input  [31:0] io_weightVec_59,
  input  [31:0] io_weightVec_60,
  input  [31:0] io_weightVec_61,
  input  [31:0] io_weightVec_62,
  input  [31:0] io_weightVec_63,
  input  [31:0] io_weightVec_64,
  input  [31:0] io_weightVec_65,
  input  [31:0] io_weightVec_66,
  input  [31:0] io_weightVec_67,
  input  [31:0] io_weightVec_68,
  input  [31:0] io_weightVec_69,
  input  [31:0] io_weightVec_70,
  input  [31:0] io_weightVec_71,
  input  [31:0] io_weightVec_72,
  input  [31:0] io_weightVec_73,
  input  [31:0] io_weightVec_74,
  input  [31:0] io_weightVec_75,
  input  [31:0] io_weightVec_76,
  input  [31:0] io_weightVec_77,
  input  [31:0] io_weightVec_78,
  input  [31:0] io_weightVec_79,
  input  [31:0] io_weightVec_80,
  input  [31:0] io_weightVec_81,
  input  [31:0] io_weightVec_82,
  input  [31:0] io_weightVec_83,
  input  [31:0] io_weightVec_84,
  input  [31:0] io_weightVec_85,
  input  [31:0] io_weightVec_86,
  input  [31:0] io_weightVec_87,
  input  [31:0] io_weightVec_88,
  input  [31:0] io_weightVec_89,
  input  [31:0] io_weightVec_90,
  input  [31:0] io_weightVec_91,
  input  [31:0] io_weightVec_92,
  input  [31:0] io_weightVec_93,
  input  [31:0] io_weightVec_94,
  input  [31:0] io_weightVec_95,
  input  [31:0] io_weightVec_96,
  input  [31:0] io_weightVec_97,
  input  [31:0] io_weightVec_98,
  input  [31:0] io_weightVec_99,
  input  [31:0] io_biasVec_0,
  input  [31:0] io_biasVec_1,
  input  [31:0] io_biasVec_2,
  input  [31:0] io_biasVec_3,
  input  [31:0] io_biasVec_4,
  input  [31:0] io_biasVec_5,
  input  [31:0] io_biasVec_6,
  input  [31:0] io_biasVec_7,
  input  [31:0] io_biasVec_8,
  input  [31:0] io_biasVec_9,
  input  [31:0] io_biasVec_10,
  input  [31:0] io_biasVec_11,
  input  [31:0] io_biasVec_12,
  input  [31:0] io_biasVec_13,
  input  [31:0] io_biasVec_14,
  input  [31:0] io_biasVec_15,
  input  [31:0] io_biasVec_16,
  input  [31:0] io_biasVec_17,
  input  [31:0] io_biasVec_18,
  input  [31:0] io_biasVec_19,
  input  [31:0] io_biasVec_20,
  input  [31:0] io_biasVec_21,
  input  [31:0] io_biasVec_22,
  input  [31:0] io_biasVec_23,
  input  [31:0] io_biasVec_24,
  input  [31:0] io_biasVec_25,
  input  [31:0] io_biasVec_26,
  input  [31:0] io_biasVec_27,
  input  [31:0] io_biasVec_28,
  input  [31:0] io_biasVec_29,
  input  [31:0] io_biasVec_30,
  input  [31:0] io_biasVec_31,
  input  [31:0] io_biasVec_32,
  input  [31:0] io_biasVec_33,
  input  [31:0] io_biasVec_34,
  input  [31:0] io_biasVec_35,
  input  [31:0] io_biasVec_36,
  input  [31:0] io_biasVec_37,
  input  [31:0] io_biasVec_38,
  input  [31:0] io_biasVec_39,
  input  [31:0] io_biasVec_40,
  input  [31:0] io_biasVec_41,
  input  [31:0] io_biasVec_42,
  input  [31:0] io_biasVec_43,
  input  [31:0] io_biasVec_44,
  input  [31:0] io_biasVec_45,
  input  [31:0] io_biasVec_46,
  input  [31:0] io_biasVec_47,
  input  [31:0] io_biasVec_48,
  input  [31:0] io_biasVec_49,
  input  [31:0] io_biasVec_50,
  input  [31:0] io_biasVec_51,
  input  [31:0] io_biasVec_52,
  input  [31:0] io_biasVec_53,
  input  [31:0] io_biasVec_54,
  input  [31:0] io_biasVec_55,
  input  [31:0] io_biasVec_56,
  input  [31:0] io_biasVec_57,
  input  [31:0] io_biasVec_58,
  input  [31:0] io_biasVec_59,
  input  [31:0] io_biasVec_60,
  input  [31:0] io_biasVec_61,
  input  [31:0] io_biasVec_62,
  input  [31:0] io_biasVec_63,
  input  [31:0] io_biasVec_64,
  input  [31:0] io_biasVec_65,
  input  [31:0] io_biasVec_66,
  input  [31:0] io_biasVec_67,
  input  [31:0] io_biasVec_68,
  input  [31:0] io_biasVec_69,
  input  [31:0] io_biasVec_70,
  input  [31:0] io_biasVec_71,
  input  [31:0] io_biasVec_72,
  input  [31:0] io_biasVec_73,
  input  [31:0] io_biasVec_74,
  input  [31:0] io_biasVec_75,
  input  [31:0] io_biasVec_76,
  input  [31:0] io_biasVec_77,
  input  [31:0] io_biasVec_78,
  input  [31:0] io_biasVec_79,
  input  [31:0] io_biasVec_80,
  input  [31:0] io_biasVec_81,
  input  [31:0] io_biasVec_82,
  input  [31:0] io_biasVec_83,
  input  [31:0] io_biasVec_84,
  input  [31:0] io_biasVec_85,
  input  [31:0] io_biasVec_86,
  input  [31:0] io_biasVec_87,
  input  [31:0] io_biasVec_88,
  input  [31:0] io_biasVec_89,
  input  [31:0] io_biasVec_90,
  input  [31:0] io_biasVec_91,
  input  [31:0] io_biasVec_92,
  input  [31:0] io_biasVec_93,
  input  [31:0] io_biasVec_94,
  input  [31:0] io_biasVec_95,
  input  [31:0] io_biasVec_96,
  input  [31:0] io_biasVec_97,
  input  [31:0] io_biasVec_98,
  input  [31:0] io_biasVec_99,
  input  [31:0] io_biasScalar,
  output [31:0] io_rawVotes
);
  wire [63:0] _T; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_2; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_3; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_5; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_6; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_8; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_9; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_11; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_12; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_13; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_14; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_15; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_16; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_18; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_19; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_21; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_22; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_24; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_25; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_26; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_27; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_28; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_29; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_31; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_32; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_34; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_35; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_37; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_38; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_39; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_40; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_41; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_42; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_44; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_45; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_47; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_48; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_50; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_51; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_52; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_53; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_54; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_55; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_57; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_58; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_60; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_61; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_63; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_64; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_65; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_66; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_67; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_68; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_70; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_71; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_73; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_74; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_76; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_77; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_78; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_79; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_80; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_81; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_83; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_84; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_86; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_87; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_89; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_90; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_91; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_92; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_93; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_94; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_96; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_97; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_99; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_100; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_102; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_103; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_104; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_105; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_106; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_107; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_109; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_110; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_112; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_113; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_115; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_116; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_117; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_118; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_119; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_120; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_122; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_123; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_125; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_126; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_128; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_129; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_130; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_131; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_132; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_133; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_135; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_136; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_138; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_139; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_141; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_142; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_143; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_144; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_145; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_146; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_148; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_149; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_151; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_152; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_154; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_155; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_156; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_157; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_158; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_159; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_161; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_162; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_164; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_165; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_167; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_168; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_169; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_170; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_171; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_172; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_174; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_175; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_177; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_178; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_180; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_181; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_182; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_183; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_184; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_185; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_187; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_188; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_190; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_191; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_193; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_194; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_195; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_196; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_197; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_198; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_200; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_201; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_203; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_204; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_206; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_207; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_208; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_209; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_210; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_211; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_213; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_214; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_216; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_217; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_219; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_220; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_221; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_222; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_223; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_224; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_226; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_227; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_229; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_230; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_232; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_233; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_234; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_235; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_236; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_237; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_239; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_240; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_242; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_243; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_245; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_246; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_247; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_248; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_249; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_250; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_252; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_253; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_255; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_256; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_258; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_259; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_260; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_261; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_262; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_263; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_265; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_266; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_268; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_269; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_271; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_272; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_273; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_274; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_275; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_276; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_278; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_279; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_281; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_282; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_284; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_285; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_286; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_287; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_288; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_289; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_291; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_292; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_294; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_295; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_297; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_298; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_299; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_300; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_301; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_302; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_304; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_305; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_307; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_308; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_310; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_311; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_312; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_313; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_314; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_315; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_317; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_318; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_320; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_321; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_323; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_324; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_325; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_326; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_327; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_328; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_330; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_331; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_333; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_334; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_336; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_337; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_338; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_339; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_340; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_341; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_343; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_344; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_346; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_347; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_349; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_350; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_351; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_352; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_353; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_354; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_356; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_357; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_359; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_360; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_362; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_363; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_364; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_365; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_366; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_367; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_369; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_370; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_372; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_373; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_375; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_376; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_377; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_378; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_379; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_380; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_382; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_383; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_385; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_386; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_388; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_389; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_390; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_391; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_392; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_393; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_395; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_396; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_398; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_399; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_401; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_402; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_403; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_404; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_405; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_406; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_408; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_409; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_411; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_412; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_414; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_415; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_416; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_417; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_418; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_419; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_421; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_422; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_424; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_425; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_427; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_428; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_429; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_430; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_431; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_432; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_434; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_435; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_437; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_438; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_440; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_441; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_442; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_443; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_444; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_445; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_447; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_448; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_450; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_451; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_453; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_454; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_455; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_456; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_457; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_458; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_460; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_461; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_463; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_464; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_466; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_467; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_468; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_469; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_470; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_471; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_473; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_474; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_476; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_477; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_479; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_480; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_481; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_482; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_483; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_484; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_486; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_487; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_489; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_490; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_492; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_493; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_494; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_495; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_496; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_497; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_499; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_500; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_502; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_503; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_505; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_506; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_507; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_508; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_509; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_510; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_512; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_513; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_515; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_516; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_518; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_519; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_520; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_521; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_522; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_523; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_525; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_526; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_528; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_529; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_531; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_532; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_533; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_534; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_535; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_536; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_538; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_539; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_541; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_542; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_544; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_545; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_546; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_547; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_548; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_549; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_551; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_552; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_554; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_555; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_557; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_558; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_559; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_560; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_561; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_562; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_564; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_565; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_567; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_568; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_570; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_571; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_572; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_573; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_574; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_575; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_577; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_578; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_580; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_581; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_583; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_584; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_585; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_586; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_587; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_588; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_590; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_591; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_593; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_594; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_596; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_597; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_598; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_599; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_600; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_601; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_603; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_604; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_606; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_607; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_609; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_610; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_611; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_612; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_613; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_614; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_616; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_617; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_619; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_620; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_622; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_623; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_624; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_625; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_626; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_627; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_629; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_630; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_632; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_633; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_635; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_636; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_637; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_638; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_639; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_640; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_642; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_643; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_645; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_646; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_648; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_649; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_650; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_651; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_652; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_653; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_655; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_656; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_658; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_659; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_661; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_662; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_663; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_664; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_665; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_666; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_668; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_669; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_671; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_672; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_674; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_675; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_676; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_677; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_678; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_679; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_681; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_682; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_684; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_685; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_687; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_688; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_689; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_690; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_691; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_692; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_694; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_695; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_697; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_698; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_700; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_701; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_702; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_703; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_704; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_705; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_707; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_708; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_710; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_711; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_713; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_714; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_715; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_716; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_717; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_718; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_720; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_721; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_723; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_724; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_726; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_727; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_728; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_729; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_730; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_731; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_733; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_734; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_736; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_737; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_739; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_740; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_741; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_742; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_743; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_744; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_746; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_747; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_749; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_750; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_752; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_753; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_754; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_755; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_756; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_757; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_759; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_760; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_762; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_763; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_765; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_766; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_767; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_768; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_769; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_770; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_772; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_773; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_775; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_776; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_778; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_779; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_780; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_781; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_782; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_783; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_785; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_786; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_788; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_789; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_791; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_792; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_793; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_794; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_795; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_796; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_798; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_799; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_801; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_802; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_804; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_805; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_806; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_807; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_808; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_809; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_811; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_812; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_814; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_815; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_817; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_818; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_819; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_820; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_821; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_822; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_824; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_825; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_827; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_828; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_830; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_831; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_832; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_833; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_834; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_835; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_837; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_838; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_840; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_841; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_843; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_844; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_845; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_846; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_847; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_848; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_850; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_851; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_853; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_854; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_856; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_857; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_858; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_859; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_860; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_861; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_863; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_864; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_866; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_867; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_869; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_870; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_871; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_872; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_873; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_874; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_876; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_877; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_879; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_880; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_882; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_883; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_884; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_885; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_886; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_887; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_889; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_890; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_892; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_893; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_895; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_896; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_897; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_898; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_899; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_900; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_902; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_903; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_905; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_906; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_908; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_909; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_910; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_911; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_912; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_913; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_915; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_916; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_918; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_919; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_921; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_922; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_923; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_924; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_925; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_926; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_928; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_929; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_931; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_932; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_934; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_935; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_936; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_937; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_938; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_939; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_941; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_942; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_944; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_945; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_947; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_948; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_949; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_950; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_951; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_952; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_954; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_955; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_957; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_958; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_960; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_961; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_962; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_963; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_964; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_965; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_967; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_968; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_970; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_971; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_973; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_974; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_975; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_976; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_977; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_978; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_980; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_981; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_983; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_984; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_986; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_987; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_988; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_989; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_990; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_991; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_993; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_994; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_996; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_997; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_999; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1000; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1001; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1002; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1003; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1004; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1006; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1007; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1009; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1010; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1012; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1013; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1014; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1015; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1016; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1017; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1019; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1020; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1022; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1023; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1025; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1026; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1027; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1028; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1029; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1030; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1032; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1033; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1035; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1036; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1038; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1039; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1040; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1041; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1042; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1043; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1045; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1046; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1048; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1049; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1051; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1052; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1053; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1054; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1055; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1056; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1058; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1059; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1061; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1062; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1064; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1065; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1066; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1067; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1068; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1069; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1071; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1072; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1074; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1075; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1077; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1078; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1079; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1080; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1081; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1082; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1084; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1085; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1087; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1088; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1090; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1091; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1092; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1093; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1094; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1095; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1097; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1098; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1100; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1101; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1103; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1104; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1105; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1106; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1107; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1108; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1110; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1111; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1113; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1114; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1116; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1117; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1118; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1119; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1120; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1121; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1123; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1124; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1126; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1127; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1129; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1130; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1131; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1132; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1133; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1134; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1136; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1137; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1139; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1140; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1142; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1143; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1144; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1145; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1146; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1147; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1149; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1150; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1152; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1153; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1155; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1156; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1157; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1158; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1159; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1160; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1162; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1163; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1165; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1166; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1168; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1169; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1170; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1171; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1172; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1173; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1175; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1176; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1178; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1179; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1181; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1182; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1183; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1184; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1185; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1186; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1188; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1189; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1191; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1192; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1194; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1195; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1196; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1197; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1198; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1199; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1201; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1202; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1204; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1205; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1207; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1208; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1209; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1210; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1211; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1212; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1214; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1215; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1217; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1218; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1220; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1221; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1222; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1223; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1224; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1225; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1227; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1228; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1230; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1231; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1233; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1234; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1235; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1236; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1237; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1238; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1240; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1241; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1243; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1244; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1246; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1247; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1248; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1249; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1250; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1251; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1253; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1254; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1256; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1257; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1259; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1260; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1261; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1262; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1263; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1264; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1266; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1267; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1269; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1270; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1272; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1273; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1274; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1275; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1276; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1277; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1279; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1280; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1282; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1283; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1285; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1286; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1287; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1288; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1289; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1290; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1292; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1293; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1295; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1296; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1298; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1299; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_2; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_3; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_0; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1301; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_0; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_4; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_5; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_1; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1304; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_1; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_6; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_7; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_2; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1307; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_2; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_8; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_9; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_3; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1310; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_3; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_10; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_11; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_4; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1313; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_4; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_12; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_13; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_5; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1316; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_5; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_14; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_15; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_6; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1319; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_6; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_16; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_17; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_7; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1322; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_7; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_18; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_19; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_8; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1325; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_8; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_20; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_21; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_9; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1328; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_9; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_22; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_23; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_10; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1331; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_10; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_24; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_25; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_11; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1334; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_11; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_26; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_27; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_12; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1337; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_12; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_28; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_29; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_13; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1340; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_13; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_30; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_31; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_14; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1343; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_14; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_32; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_33; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_15; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1346; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_15; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_34; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_35; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_16; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1349; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_16; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_36; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_37; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_17; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1352; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_17; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_38; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_39; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_18; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1355; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_18; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_40; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_41; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_19; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1358; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_19; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_42; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_43; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_20; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1361; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_20; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_44; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_45; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_21; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1364; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_21; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_46; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_47; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_22; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1367; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_22; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_48; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_49; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_23; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1370; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_23; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_50; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_51; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_24; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1373; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_24; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_52; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_53; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_25; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1376; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_25; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_54; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_55; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_26; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1379; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_26; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_56; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_57; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_27; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1382; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_27; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_58; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_59; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_28; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1385; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_28; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_60; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_61; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_29; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1388; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_29; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_62; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_63; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_30; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1391; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_30; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_64; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_65; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_31; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1394; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_31; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_66; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_67; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_32; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1397; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_32; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_68; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_69; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_33; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1400; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_33; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_70; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_71; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_34; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1403; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_34; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_72; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_73; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_35; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1406; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_35; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_74; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_75; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_36; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1409; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_36; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_76; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_77; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_37; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1412; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_37; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_78; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_79; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_38; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1415; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_38; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_80; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_81; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_39; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1418; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_39; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_82; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_83; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_40; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1421; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_40; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_84; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_85; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_41; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1424; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_41; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_86; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_87; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_42; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1427; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_42; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_88; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_89; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_43; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1430; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_43; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_90; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_91; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_44; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1433; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_44; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_92; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_93; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_45; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1436; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_45; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_94; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_95; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_46; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1439; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_46; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_96; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_97; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_47; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1442; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_47; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_98; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_99; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_48; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1445; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_48; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_100; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_101; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_49; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1448; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_49; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_102; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_103; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_50; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1451; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_50; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_104; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_105; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_51; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1454; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_51; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_106; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_107; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_52; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1457; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_52; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_108; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_109; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_53; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1460; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_53; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_110; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_111; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_54; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1463; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_54; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_112; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_113; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_55; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1466; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_55; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_114; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_115; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_56; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1469; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_56; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_116; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_117; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_57; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1472; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_57; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_118; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_119; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_58; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1475; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_58; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_120; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_121; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_59; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1478; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_59; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_122; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_123; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_60; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1481; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_60; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_124; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_125; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_61; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1484; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_61; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_126; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_127; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_62; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1487; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_62; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_128; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_129; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_63; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1490; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_63; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_130; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_131; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_64; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1493; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_64; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_132; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_133; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_65; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1496; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_65; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_134; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_135; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_66; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1499; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_66; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_136; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_137; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_67; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1502; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_67; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_138; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_139; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_68; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1505; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_68; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_140; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_141; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_69; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1508; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_69; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_142; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_143; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_70; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1511; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_70; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_144; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_145; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_71; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1514; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_71; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_146; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_147; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_72; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1517; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_72; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_148; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_149; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_73; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1520; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_73; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_150; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_151; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_74; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1523; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_74; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_152; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_153; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_75; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1526; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_75; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_154; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_155; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_76; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1529; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_76; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_156; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_157; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_77; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1532; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_77; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_158; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_159; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_78; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1535; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_78; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_160; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_161; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_79; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1538; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_79; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_162; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_163; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_80; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1541; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_80; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_164; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_165; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_81; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1544; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_81; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_166; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_167; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_82; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1547; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_82; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_168; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_169; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_83; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1550; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_83; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_170; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_171; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_84; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1553; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_84; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_172; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_173; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_85; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1556; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_85; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_174; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_175; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_86; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1559; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_86; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_176; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_177; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_87; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1562; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_87; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_178; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_179; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_88; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1565; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_88; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_180; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_181; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_89; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1568; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_89; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_182; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_183; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_90; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1571; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_90; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_184; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_185; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_91; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1574; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_91; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_186; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_187; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_92; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1577; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_92; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_188; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_189; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_93; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1580; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_93; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_190; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_191; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_94; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1583; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_94; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_192; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_193; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_95; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1586; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_95; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_194; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_195; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_96; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1589; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_96; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_196; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_197; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_97; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1592; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_97; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_198; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_199; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_98; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1595; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_98; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_200; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _GEN_201; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] inputWeighted_99; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  wire [31:0] _T_1598; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] biased_99; // @[FixedPointTypeClass.scala 21:58]
  wire  _T_1600; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_0; // @[neuralNet.scala 62:26]
  wire  _T_1602; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_1; // @[neuralNet.scala 62:26]
  wire  _T_1604; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_2; // @[neuralNet.scala 62:26]
  wire  _T_1606; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_3; // @[neuralNet.scala 62:26]
  wire  _T_1608; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_4; // @[neuralNet.scala 62:26]
  wire  _T_1610; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_5; // @[neuralNet.scala 62:26]
  wire  _T_1612; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_6; // @[neuralNet.scala 62:26]
  wire  _T_1614; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_7; // @[neuralNet.scala 62:26]
  wire  _T_1616; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_8; // @[neuralNet.scala 62:26]
  wire  _T_1618; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_9; // @[neuralNet.scala 62:26]
  wire  _T_1620; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_10; // @[neuralNet.scala 62:26]
  wire  _T_1622; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_11; // @[neuralNet.scala 62:26]
  wire  _T_1624; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_12; // @[neuralNet.scala 62:26]
  wire  _T_1626; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_13; // @[neuralNet.scala 62:26]
  wire  _T_1628; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_14; // @[neuralNet.scala 62:26]
  wire  _T_1630; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_15; // @[neuralNet.scala 62:26]
  wire  _T_1632; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_16; // @[neuralNet.scala 62:26]
  wire  _T_1634; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_17; // @[neuralNet.scala 62:26]
  wire  _T_1636; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_18; // @[neuralNet.scala 62:26]
  wire  _T_1638; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_19; // @[neuralNet.scala 62:26]
  wire  _T_1640; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_20; // @[neuralNet.scala 62:26]
  wire  _T_1642; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_21; // @[neuralNet.scala 62:26]
  wire  _T_1644; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_22; // @[neuralNet.scala 62:26]
  wire  _T_1646; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_23; // @[neuralNet.scala 62:26]
  wire  _T_1648; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_24; // @[neuralNet.scala 62:26]
  wire  _T_1650; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_25; // @[neuralNet.scala 62:26]
  wire  _T_1652; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_26; // @[neuralNet.scala 62:26]
  wire  _T_1654; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_27; // @[neuralNet.scala 62:26]
  wire  _T_1656; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_28; // @[neuralNet.scala 62:26]
  wire  _T_1658; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_29; // @[neuralNet.scala 62:26]
  wire  _T_1660; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_30; // @[neuralNet.scala 62:26]
  wire  _T_1662; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_31; // @[neuralNet.scala 62:26]
  wire  _T_1664; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_32; // @[neuralNet.scala 62:26]
  wire  _T_1666; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_33; // @[neuralNet.scala 62:26]
  wire  _T_1668; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_34; // @[neuralNet.scala 62:26]
  wire  _T_1670; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_35; // @[neuralNet.scala 62:26]
  wire  _T_1672; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_36; // @[neuralNet.scala 62:26]
  wire  _T_1674; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_37; // @[neuralNet.scala 62:26]
  wire  _T_1676; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_38; // @[neuralNet.scala 62:26]
  wire  _T_1678; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_39; // @[neuralNet.scala 62:26]
  wire  _T_1680; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_40; // @[neuralNet.scala 62:26]
  wire  _T_1682; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_41; // @[neuralNet.scala 62:26]
  wire  _T_1684; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_42; // @[neuralNet.scala 62:26]
  wire  _T_1686; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_43; // @[neuralNet.scala 62:26]
  wire  _T_1688; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_44; // @[neuralNet.scala 62:26]
  wire  _T_1690; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_45; // @[neuralNet.scala 62:26]
  wire  _T_1692; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_46; // @[neuralNet.scala 62:26]
  wire  _T_1694; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_47; // @[neuralNet.scala 62:26]
  wire  _T_1696; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_48; // @[neuralNet.scala 62:26]
  wire  _T_1698; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_49; // @[neuralNet.scala 62:26]
  wire  _T_1700; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_50; // @[neuralNet.scala 62:26]
  wire  _T_1702; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_51; // @[neuralNet.scala 62:26]
  wire  _T_1704; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_52; // @[neuralNet.scala 62:26]
  wire  _T_1706; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_53; // @[neuralNet.scala 62:26]
  wire  _T_1708; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_54; // @[neuralNet.scala 62:26]
  wire  _T_1710; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_55; // @[neuralNet.scala 62:26]
  wire  _T_1712; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_56; // @[neuralNet.scala 62:26]
  wire  _T_1714; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_57; // @[neuralNet.scala 62:26]
  wire  _T_1716; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_58; // @[neuralNet.scala 62:26]
  wire  _T_1718; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_59; // @[neuralNet.scala 62:26]
  wire  _T_1720; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_60; // @[neuralNet.scala 62:26]
  wire  _T_1722; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_61; // @[neuralNet.scala 62:26]
  wire  _T_1724; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_62; // @[neuralNet.scala 62:26]
  wire  _T_1726; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_63; // @[neuralNet.scala 62:26]
  wire  _T_1728; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_64; // @[neuralNet.scala 62:26]
  wire  _T_1730; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_65; // @[neuralNet.scala 62:26]
  wire  _T_1732; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_66; // @[neuralNet.scala 62:26]
  wire  _T_1734; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_67; // @[neuralNet.scala 62:26]
  wire  _T_1736; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_68; // @[neuralNet.scala 62:26]
  wire  _T_1738; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_69; // @[neuralNet.scala 62:26]
  wire  _T_1740; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_70; // @[neuralNet.scala 62:26]
  wire  _T_1742; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_71; // @[neuralNet.scala 62:26]
  wire  _T_1744; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_72; // @[neuralNet.scala 62:26]
  wire  _T_1746; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_73; // @[neuralNet.scala 62:26]
  wire  _T_1748; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_74; // @[neuralNet.scala 62:26]
  wire  _T_1750; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_75; // @[neuralNet.scala 62:26]
  wire  _T_1752; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_76; // @[neuralNet.scala 62:26]
  wire  _T_1754; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_77; // @[neuralNet.scala 62:26]
  wire  _T_1756; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_78; // @[neuralNet.scala 62:26]
  wire  _T_1758; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_79; // @[neuralNet.scala 62:26]
  wire  _T_1760; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_80; // @[neuralNet.scala 62:26]
  wire  _T_1762; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_81; // @[neuralNet.scala 62:26]
  wire  _T_1764; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_82; // @[neuralNet.scala 62:26]
  wire  _T_1766; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_83; // @[neuralNet.scala 62:26]
  wire  _T_1768; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_84; // @[neuralNet.scala 62:26]
  wire  _T_1770; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_85; // @[neuralNet.scala 62:26]
  wire  _T_1772; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_86; // @[neuralNet.scala 62:26]
  wire  _T_1774; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_87; // @[neuralNet.scala 62:26]
  wire  _T_1776; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_88; // @[neuralNet.scala 62:26]
  wire  _T_1778; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_89; // @[neuralNet.scala 62:26]
  wire  _T_1780; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_90; // @[neuralNet.scala 62:26]
  wire  _T_1782; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_91; // @[neuralNet.scala 62:26]
  wire  _T_1784; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_92; // @[neuralNet.scala 62:26]
  wire  _T_1786; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_93; // @[neuralNet.scala 62:26]
  wire  _T_1788; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_94; // @[neuralNet.scala 62:26]
  wire  _T_1790; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_95; // @[neuralNet.scala 62:26]
  wire  _T_1792; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_96; // @[neuralNet.scala 62:26]
  wire  _T_1794; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_97; // @[neuralNet.scala 62:26]
  wire  _T_1796; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_98; // @[neuralNet.scala 62:26]
  wire  _T_1798; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] hiddenLayer_99; // @[neuralNet.scala 62:26]
  wire [63:0] _T_1800; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1801; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1802; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1803; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1804; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1805; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1806; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1807; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1808; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1809; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1810; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1811; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1812; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1813; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1814; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1815; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1816; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1817; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1818; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1819; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1820; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1821; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1822; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1823; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1824; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1825; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1826; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1827; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1828; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1829; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1830; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1831; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1832; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1833; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1834; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1835; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1836; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1837; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1838; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1839; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1840; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1841; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1842; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1843; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1844; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1845; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1846; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1847; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1848; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1849; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1850; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1851; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1852; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1853; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1854; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1855; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1856; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1857; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1858; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1859; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1860; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1861; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1862; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1863; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1864; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1865; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1866; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1867; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1868; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1869; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1870; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1871; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1872; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1873; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1874; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1875; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1876; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1877; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1878; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1879; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1880; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1881; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1882; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1883; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1884; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1885; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1886; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1887; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1888; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1889; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1890; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1891; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1892; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1893; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1894; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1895; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1896; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1897; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1898; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1899; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1901; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1902; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1904; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1905; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1907; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1908; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1910; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1911; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1913; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1914; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1916; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1917; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1919; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1920; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1922; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1923; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1925; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1926; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1928; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1929; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1931; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1932; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1934; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1935; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1937; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1938; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1940; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1941; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1943; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1944; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1946; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1947; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1949; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1950; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1952; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1953; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1955; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1956; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1958; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1959; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1961; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1962; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1964; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1965; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1967; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1968; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1970; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1971; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1973; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1974; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1976; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1977; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1979; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1980; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1982; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1983; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1985; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1986; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1988; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1989; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1991; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1992; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1994; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1995; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1997; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1998; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2000; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2001; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2003; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2004; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2006; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2007; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2009; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2010; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2012; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2013; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2015; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2016; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2018; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2019; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2021; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2022; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2024; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2025; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2027; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2028; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2030; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2031; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2033; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2034; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2036; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2037; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2039; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2040; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2042; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2043; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2045; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2046; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2048; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2049; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2051; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2052; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2054; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2055; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2057; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2058; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2060; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2061; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2063; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2064; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2066; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2067; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2069; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2070; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2072; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2073; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2075; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2076; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2078; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2079; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2081; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2082; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2084; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2085; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2087; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2088; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2090; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2091; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2093; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2094; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2096; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2097; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2099; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2100; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2102; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2103; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2105; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2106; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2108; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2109; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2111; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2112; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2114; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2115; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2117; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2118; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2120; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2121; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2123; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2124; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2126; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2127; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2129; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2130; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2132; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2133; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2135; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2136; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2138; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2139; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2141; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2142; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2144; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2145; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2147; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2148; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2150; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2151; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2153; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2154; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2156; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2157; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2159; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2160; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2162; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2163; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2165; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2166; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2168; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2169; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2171; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2172; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2174; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2175; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2177; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2178; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2180; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2181; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2183; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2184; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2186; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2187; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2189; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2190; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2192; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2193; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2195; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_2196; // @[FixedPointTypeClass.scala 21:58]
  wire [55:0] _GEN_202; // @[neuralNet.scala 66:24 neuralNet.scala 68:16 neuralNet.scala 68:16 neuralNet.scala 68:16 neuralNet.scala 68:16]
  wire [31:0] _GEN_203; // @[neuralNet.scala 66:24 neuralNet.scala 68:16 neuralNet.scala 68:16 neuralNet.scala 68:16 neuralNet.scala 68:16]
  wire [31:0] dotProduct; // @[neuralNet.scala 66:24 neuralNet.scala 68:16 neuralNet.scala 68:16 neuralNet.scala 68:16 neuralNet.scala 68:16]
  wire [31:0] _T_3389; // @[FixedPointTypeClass.scala 21:58]
  wire [31:0] actualPreReLU; // @[FixedPointTypeClass.scala 21:58]
  wire  _T_3391; // @[FixedPointTypeClass.scala 56:59]
  wire [31:0] actualVotes; // @[neuralNet.scala 75:21]
  wire  finalPredict; // @[FixedPointTypeClass.scala 56:59]
  reg [31:0] rawVotesReg; // @[Reg.scala 11:16]
  reg [31:0] _RAND_0;
  reg  outReg; // @[Reg.scala 11:16]
  reg [31:0] _RAND_1;
  reg  valReg; // @[neuralNet.scala 83:23]
  reg [31:0] _RAND_2;
  assign _T = $signed(io_in_bits_0) * $signed(io_weightMatrix_0_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1 = $signed(io_in_bits_1) * $signed(io_weightMatrix_0_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_2 = $signed(io_in_bits_2) * $signed(io_weightMatrix_0_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_3 = $signed(io_in_bits_3) * $signed(io_weightMatrix_0_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_5 = $signed(_T) + $signed(_T_1); // @[FixedPointTypeClass.scala 21:58]
  assign _T_6 = $signed(_T_5); // @[FixedPointTypeClass.scala 21:58]
  assign _T_8 = $signed(_T_6) + $signed(_T_2); // @[FixedPointTypeClass.scala 21:58]
  assign _T_9 = $signed(_T_8); // @[FixedPointTypeClass.scala 21:58]
  assign _T_11 = $signed(_T_9) + $signed(_T_3); // @[FixedPointTypeClass.scala 21:58]
  assign _T_12 = $signed(_T_11); // @[FixedPointTypeClass.scala 21:58]
  assign _T_13 = $signed(io_in_bits_0) * $signed(io_weightMatrix_1_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_14 = $signed(io_in_bits_1) * $signed(io_weightMatrix_1_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_15 = $signed(io_in_bits_2) * $signed(io_weightMatrix_1_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_16 = $signed(io_in_bits_3) * $signed(io_weightMatrix_1_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_18 = $signed(_T_13) + $signed(_T_14); // @[FixedPointTypeClass.scala 21:58]
  assign _T_19 = $signed(_T_18); // @[FixedPointTypeClass.scala 21:58]
  assign _T_21 = $signed(_T_19) + $signed(_T_15); // @[FixedPointTypeClass.scala 21:58]
  assign _T_22 = $signed(_T_21); // @[FixedPointTypeClass.scala 21:58]
  assign _T_24 = $signed(_T_22) + $signed(_T_16); // @[FixedPointTypeClass.scala 21:58]
  assign _T_25 = $signed(_T_24); // @[FixedPointTypeClass.scala 21:58]
  assign _T_26 = $signed(io_in_bits_0) * $signed(io_weightMatrix_2_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_27 = $signed(io_in_bits_1) * $signed(io_weightMatrix_2_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_28 = $signed(io_in_bits_2) * $signed(io_weightMatrix_2_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_29 = $signed(io_in_bits_3) * $signed(io_weightMatrix_2_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_31 = $signed(_T_26) + $signed(_T_27); // @[FixedPointTypeClass.scala 21:58]
  assign _T_32 = $signed(_T_31); // @[FixedPointTypeClass.scala 21:58]
  assign _T_34 = $signed(_T_32) + $signed(_T_28); // @[FixedPointTypeClass.scala 21:58]
  assign _T_35 = $signed(_T_34); // @[FixedPointTypeClass.scala 21:58]
  assign _T_37 = $signed(_T_35) + $signed(_T_29); // @[FixedPointTypeClass.scala 21:58]
  assign _T_38 = $signed(_T_37); // @[FixedPointTypeClass.scala 21:58]
  assign _T_39 = $signed(io_in_bits_0) * $signed(io_weightMatrix_3_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_40 = $signed(io_in_bits_1) * $signed(io_weightMatrix_3_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_41 = $signed(io_in_bits_2) * $signed(io_weightMatrix_3_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_42 = $signed(io_in_bits_3) * $signed(io_weightMatrix_3_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_44 = $signed(_T_39) + $signed(_T_40); // @[FixedPointTypeClass.scala 21:58]
  assign _T_45 = $signed(_T_44); // @[FixedPointTypeClass.scala 21:58]
  assign _T_47 = $signed(_T_45) + $signed(_T_41); // @[FixedPointTypeClass.scala 21:58]
  assign _T_48 = $signed(_T_47); // @[FixedPointTypeClass.scala 21:58]
  assign _T_50 = $signed(_T_48) + $signed(_T_42); // @[FixedPointTypeClass.scala 21:58]
  assign _T_51 = $signed(_T_50); // @[FixedPointTypeClass.scala 21:58]
  assign _T_52 = $signed(io_in_bits_0) * $signed(io_weightMatrix_4_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_53 = $signed(io_in_bits_1) * $signed(io_weightMatrix_4_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_54 = $signed(io_in_bits_2) * $signed(io_weightMatrix_4_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_55 = $signed(io_in_bits_3) * $signed(io_weightMatrix_4_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_57 = $signed(_T_52) + $signed(_T_53); // @[FixedPointTypeClass.scala 21:58]
  assign _T_58 = $signed(_T_57); // @[FixedPointTypeClass.scala 21:58]
  assign _T_60 = $signed(_T_58) + $signed(_T_54); // @[FixedPointTypeClass.scala 21:58]
  assign _T_61 = $signed(_T_60); // @[FixedPointTypeClass.scala 21:58]
  assign _T_63 = $signed(_T_61) + $signed(_T_55); // @[FixedPointTypeClass.scala 21:58]
  assign _T_64 = $signed(_T_63); // @[FixedPointTypeClass.scala 21:58]
  assign _T_65 = $signed(io_in_bits_0) * $signed(io_weightMatrix_5_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_66 = $signed(io_in_bits_1) * $signed(io_weightMatrix_5_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_67 = $signed(io_in_bits_2) * $signed(io_weightMatrix_5_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_68 = $signed(io_in_bits_3) * $signed(io_weightMatrix_5_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_70 = $signed(_T_65) + $signed(_T_66); // @[FixedPointTypeClass.scala 21:58]
  assign _T_71 = $signed(_T_70); // @[FixedPointTypeClass.scala 21:58]
  assign _T_73 = $signed(_T_71) + $signed(_T_67); // @[FixedPointTypeClass.scala 21:58]
  assign _T_74 = $signed(_T_73); // @[FixedPointTypeClass.scala 21:58]
  assign _T_76 = $signed(_T_74) + $signed(_T_68); // @[FixedPointTypeClass.scala 21:58]
  assign _T_77 = $signed(_T_76); // @[FixedPointTypeClass.scala 21:58]
  assign _T_78 = $signed(io_in_bits_0) * $signed(io_weightMatrix_6_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_79 = $signed(io_in_bits_1) * $signed(io_weightMatrix_6_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_80 = $signed(io_in_bits_2) * $signed(io_weightMatrix_6_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_81 = $signed(io_in_bits_3) * $signed(io_weightMatrix_6_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_83 = $signed(_T_78) + $signed(_T_79); // @[FixedPointTypeClass.scala 21:58]
  assign _T_84 = $signed(_T_83); // @[FixedPointTypeClass.scala 21:58]
  assign _T_86 = $signed(_T_84) + $signed(_T_80); // @[FixedPointTypeClass.scala 21:58]
  assign _T_87 = $signed(_T_86); // @[FixedPointTypeClass.scala 21:58]
  assign _T_89 = $signed(_T_87) + $signed(_T_81); // @[FixedPointTypeClass.scala 21:58]
  assign _T_90 = $signed(_T_89); // @[FixedPointTypeClass.scala 21:58]
  assign _T_91 = $signed(io_in_bits_0) * $signed(io_weightMatrix_7_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_92 = $signed(io_in_bits_1) * $signed(io_weightMatrix_7_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_93 = $signed(io_in_bits_2) * $signed(io_weightMatrix_7_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_94 = $signed(io_in_bits_3) * $signed(io_weightMatrix_7_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_96 = $signed(_T_91) + $signed(_T_92); // @[FixedPointTypeClass.scala 21:58]
  assign _T_97 = $signed(_T_96); // @[FixedPointTypeClass.scala 21:58]
  assign _T_99 = $signed(_T_97) + $signed(_T_93); // @[FixedPointTypeClass.scala 21:58]
  assign _T_100 = $signed(_T_99); // @[FixedPointTypeClass.scala 21:58]
  assign _T_102 = $signed(_T_100) + $signed(_T_94); // @[FixedPointTypeClass.scala 21:58]
  assign _T_103 = $signed(_T_102); // @[FixedPointTypeClass.scala 21:58]
  assign _T_104 = $signed(io_in_bits_0) * $signed(io_weightMatrix_8_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_105 = $signed(io_in_bits_1) * $signed(io_weightMatrix_8_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_106 = $signed(io_in_bits_2) * $signed(io_weightMatrix_8_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_107 = $signed(io_in_bits_3) * $signed(io_weightMatrix_8_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_109 = $signed(_T_104) + $signed(_T_105); // @[FixedPointTypeClass.scala 21:58]
  assign _T_110 = $signed(_T_109); // @[FixedPointTypeClass.scala 21:58]
  assign _T_112 = $signed(_T_110) + $signed(_T_106); // @[FixedPointTypeClass.scala 21:58]
  assign _T_113 = $signed(_T_112); // @[FixedPointTypeClass.scala 21:58]
  assign _T_115 = $signed(_T_113) + $signed(_T_107); // @[FixedPointTypeClass.scala 21:58]
  assign _T_116 = $signed(_T_115); // @[FixedPointTypeClass.scala 21:58]
  assign _T_117 = $signed(io_in_bits_0) * $signed(io_weightMatrix_9_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_118 = $signed(io_in_bits_1) * $signed(io_weightMatrix_9_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_119 = $signed(io_in_bits_2) * $signed(io_weightMatrix_9_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_120 = $signed(io_in_bits_3) * $signed(io_weightMatrix_9_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_122 = $signed(_T_117) + $signed(_T_118); // @[FixedPointTypeClass.scala 21:58]
  assign _T_123 = $signed(_T_122); // @[FixedPointTypeClass.scala 21:58]
  assign _T_125 = $signed(_T_123) + $signed(_T_119); // @[FixedPointTypeClass.scala 21:58]
  assign _T_126 = $signed(_T_125); // @[FixedPointTypeClass.scala 21:58]
  assign _T_128 = $signed(_T_126) + $signed(_T_120); // @[FixedPointTypeClass.scala 21:58]
  assign _T_129 = $signed(_T_128); // @[FixedPointTypeClass.scala 21:58]
  assign _T_130 = $signed(io_in_bits_0) * $signed(io_weightMatrix_10_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_131 = $signed(io_in_bits_1) * $signed(io_weightMatrix_10_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_132 = $signed(io_in_bits_2) * $signed(io_weightMatrix_10_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_133 = $signed(io_in_bits_3) * $signed(io_weightMatrix_10_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_135 = $signed(_T_130) + $signed(_T_131); // @[FixedPointTypeClass.scala 21:58]
  assign _T_136 = $signed(_T_135); // @[FixedPointTypeClass.scala 21:58]
  assign _T_138 = $signed(_T_136) + $signed(_T_132); // @[FixedPointTypeClass.scala 21:58]
  assign _T_139 = $signed(_T_138); // @[FixedPointTypeClass.scala 21:58]
  assign _T_141 = $signed(_T_139) + $signed(_T_133); // @[FixedPointTypeClass.scala 21:58]
  assign _T_142 = $signed(_T_141); // @[FixedPointTypeClass.scala 21:58]
  assign _T_143 = $signed(io_in_bits_0) * $signed(io_weightMatrix_11_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_144 = $signed(io_in_bits_1) * $signed(io_weightMatrix_11_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_145 = $signed(io_in_bits_2) * $signed(io_weightMatrix_11_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_146 = $signed(io_in_bits_3) * $signed(io_weightMatrix_11_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_148 = $signed(_T_143) + $signed(_T_144); // @[FixedPointTypeClass.scala 21:58]
  assign _T_149 = $signed(_T_148); // @[FixedPointTypeClass.scala 21:58]
  assign _T_151 = $signed(_T_149) + $signed(_T_145); // @[FixedPointTypeClass.scala 21:58]
  assign _T_152 = $signed(_T_151); // @[FixedPointTypeClass.scala 21:58]
  assign _T_154 = $signed(_T_152) + $signed(_T_146); // @[FixedPointTypeClass.scala 21:58]
  assign _T_155 = $signed(_T_154); // @[FixedPointTypeClass.scala 21:58]
  assign _T_156 = $signed(io_in_bits_0) * $signed(io_weightMatrix_12_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_157 = $signed(io_in_bits_1) * $signed(io_weightMatrix_12_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_158 = $signed(io_in_bits_2) * $signed(io_weightMatrix_12_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_159 = $signed(io_in_bits_3) * $signed(io_weightMatrix_12_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_161 = $signed(_T_156) + $signed(_T_157); // @[FixedPointTypeClass.scala 21:58]
  assign _T_162 = $signed(_T_161); // @[FixedPointTypeClass.scala 21:58]
  assign _T_164 = $signed(_T_162) + $signed(_T_158); // @[FixedPointTypeClass.scala 21:58]
  assign _T_165 = $signed(_T_164); // @[FixedPointTypeClass.scala 21:58]
  assign _T_167 = $signed(_T_165) + $signed(_T_159); // @[FixedPointTypeClass.scala 21:58]
  assign _T_168 = $signed(_T_167); // @[FixedPointTypeClass.scala 21:58]
  assign _T_169 = $signed(io_in_bits_0) * $signed(io_weightMatrix_13_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_170 = $signed(io_in_bits_1) * $signed(io_weightMatrix_13_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_171 = $signed(io_in_bits_2) * $signed(io_weightMatrix_13_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_172 = $signed(io_in_bits_3) * $signed(io_weightMatrix_13_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_174 = $signed(_T_169) + $signed(_T_170); // @[FixedPointTypeClass.scala 21:58]
  assign _T_175 = $signed(_T_174); // @[FixedPointTypeClass.scala 21:58]
  assign _T_177 = $signed(_T_175) + $signed(_T_171); // @[FixedPointTypeClass.scala 21:58]
  assign _T_178 = $signed(_T_177); // @[FixedPointTypeClass.scala 21:58]
  assign _T_180 = $signed(_T_178) + $signed(_T_172); // @[FixedPointTypeClass.scala 21:58]
  assign _T_181 = $signed(_T_180); // @[FixedPointTypeClass.scala 21:58]
  assign _T_182 = $signed(io_in_bits_0) * $signed(io_weightMatrix_14_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_183 = $signed(io_in_bits_1) * $signed(io_weightMatrix_14_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_184 = $signed(io_in_bits_2) * $signed(io_weightMatrix_14_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_185 = $signed(io_in_bits_3) * $signed(io_weightMatrix_14_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_187 = $signed(_T_182) + $signed(_T_183); // @[FixedPointTypeClass.scala 21:58]
  assign _T_188 = $signed(_T_187); // @[FixedPointTypeClass.scala 21:58]
  assign _T_190 = $signed(_T_188) + $signed(_T_184); // @[FixedPointTypeClass.scala 21:58]
  assign _T_191 = $signed(_T_190); // @[FixedPointTypeClass.scala 21:58]
  assign _T_193 = $signed(_T_191) + $signed(_T_185); // @[FixedPointTypeClass.scala 21:58]
  assign _T_194 = $signed(_T_193); // @[FixedPointTypeClass.scala 21:58]
  assign _T_195 = $signed(io_in_bits_0) * $signed(io_weightMatrix_15_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_196 = $signed(io_in_bits_1) * $signed(io_weightMatrix_15_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_197 = $signed(io_in_bits_2) * $signed(io_weightMatrix_15_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_198 = $signed(io_in_bits_3) * $signed(io_weightMatrix_15_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_200 = $signed(_T_195) + $signed(_T_196); // @[FixedPointTypeClass.scala 21:58]
  assign _T_201 = $signed(_T_200); // @[FixedPointTypeClass.scala 21:58]
  assign _T_203 = $signed(_T_201) + $signed(_T_197); // @[FixedPointTypeClass.scala 21:58]
  assign _T_204 = $signed(_T_203); // @[FixedPointTypeClass.scala 21:58]
  assign _T_206 = $signed(_T_204) + $signed(_T_198); // @[FixedPointTypeClass.scala 21:58]
  assign _T_207 = $signed(_T_206); // @[FixedPointTypeClass.scala 21:58]
  assign _T_208 = $signed(io_in_bits_0) * $signed(io_weightMatrix_16_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_209 = $signed(io_in_bits_1) * $signed(io_weightMatrix_16_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_210 = $signed(io_in_bits_2) * $signed(io_weightMatrix_16_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_211 = $signed(io_in_bits_3) * $signed(io_weightMatrix_16_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_213 = $signed(_T_208) + $signed(_T_209); // @[FixedPointTypeClass.scala 21:58]
  assign _T_214 = $signed(_T_213); // @[FixedPointTypeClass.scala 21:58]
  assign _T_216 = $signed(_T_214) + $signed(_T_210); // @[FixedPointTypeClass.scala 21:58]
  assign _T_217 = $signed(_T_216); // @[FixedPointTypeClass.scala 21:58]
  assign _T_219 = $signed(_T_217) + $signed(_T_211); // @[FixedPointTypeClass.scala 21:58]
  assign _T_220 = $signed(_T_219); // @[FixedPointTypeClass.scala 21:58]
  assign _T_221 = $signed(io_in_bits_0) * $signed(io_weightMatrix_17_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_222 = $signed(io_in_bits_1) * $signed(io_weightMatrix_17_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_223 = $signed(io_in_bits_2) * $signed(io_weightMatrix_17_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_224 = $signed(io_in_bits_3) * $signed(io_weightMatrix_17_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_226 = $signed(_T_221) + $signed(_T_222); // @[FixedPointTypeClass.scala 21:58]
  assign _T_227 = $signed(_T_226); // @[FixedPointTypeClass.scala 21:58]
  assign _T_229 = $signed(_T_227) + $signed(_T_223); // @[FixedPointTypeClass.scala 21:58]
  assign _T_230 = $signed(_T_229); // @[FixedPointTypeClass.scala 21:58]
  assign _T_232 = $signed(_T_230) + $signed(_T_224); // @[FixedPointTypeClass.scala 21:58]
  assign _T_233 = $signed(_T_232); // @[FixedPointTypeClass.scala 21:58]
  assign _T_234 = $signed(io_in_bits_0) * $signed(io_weightMatrix_18_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_235 = $signed(io_in_bits_1) * $signed(io_weightMatrix_18_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_236 = $signed(io_in_bits_2) * $signed(io_weightMatrix_18_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_237 = $signed(io_in_bits_3) * $signed(io_weightMatrix_18_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_239 = $signed(_T_234) + $signed(_T_235); // @[FixedPointTypeClass.scala 21:58]
  assign _T_240 = $signed(_T_239); // @[FixedPointTypeClass.scala 21:58]
  assign _T_242 = $signed(_T_240) + $signed(_T_236); // @[FixedPointTypeClass.scala 21:58]
  assign _T_243 = $signed(_T_242); // @[FixedPointTypeClass.scala 21:58]
  assign _T_245 = $signed(_T_243) + $signed(_T_237); // @[FixedPointTypeClass.scala 21:58]
  assign _T_246 = $signed(_T_245); // @[FixedPointTypeClass.scala 21:58]
  assign _T_247 = $signed(io_in_bits_0) * $signed(io_weightMatrix_19_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_248 = $signed(io_in_bits_1) * $signed(io_weightMatrix_19_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_249 = $signed(io_in_bits_2) * $signed(io_weightMatrix_19_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_250 = $signed(io_in_bits_3) * $signed(io_weightMatrix_19_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_252 = $signed(_T_247) + $signed(_T_248); // @[FixedPointTypeClass.scala 21:58]
  assign _T_253 = $signed(_T_252); // @[FixedPointTypeClass.scala 21:58]
  assign _T_255 = $signed(_T_253) + $signed(_T_249); // @[FixedPointTypeClass.scala 21:58]
  assign _T_256 = $signed(_T_255); // @[FixedPointTypeClass.scala 21:58]
  assign _T_258 = $signed(_T_256) + $signed(_T_250); // @[FixedPointTypeClass.scala 21:58]
  assign _T_259 = $signed(_T_258); // @[FixedPointTypeClass.scala 21:58]
  assign _T_260 = $signed(io_in_bits_0) * $signed(io_weightMatrix_20_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_261 = $signed(io_in_bits_1) * $signed(io_weightMatrix_20_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_262 = $signed(io_in_bits_2) * $signed(io_weightMatrix_20_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_263 = $signed(io_in_bits_3) * $signed(io_weightMatrix_20_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_265 = $signed(_T_260) + $signed(_T_261); // @[FixedPointTypeClass.scala 21:58]
  assign _T_266 = $signed(_T_265); // @[FixedPointTypeClass.scala 21:58]
  assign _T_268 = $signed(_T_266) + $signed(_T_262); // @[FixedPointTypeClass.scala 21:58]
  assign _T_269 = $signed(_T_268); // @[FixedPointTypeClass.scala 21:58]
  assign _T_271 = $signed(_T_269) + $signed(_T_263); // @[FixedPointTypeClass.scala 21:58]
  assign _T_272 = $signed(_T_271); // @[FixedPointTypeClass.scala 21:58]
  assign _T_273 = $signed(io_in_bits_0) * $signed(io_weightMatrix_21_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_274 = $signed(io_in_bits_1) * $signed(io_weightMatrix_21_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_275 = $signed(io_in_bits_2) * $signed(io_weightMatrix_21_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_276 = $signed(io_in_bits_3) * $signed(io_weightMatrix_21_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_278 = $signed(_T_273) + $signed(_T_274); // @[FixedPointTypeClass.scala 21:58]
  assign _T_279 = $signed(_T_278); // @[FixedPointTypeClass.scala 21:58]
  assign _T_281 = $signed(_T_279) + $signed(_T_275); // @[FixedPointTypeClass.scala 21:58]
  assign _T_282 = $signed(_T_281); // @[FixedPointTypeClass.scala 21:58]
  assign _T_284 = $signed(_T_282) + $signed(_T_276); // @[FixedPointTypeClass.scala 21:58]
  assign _T_285 = $signed(_T_284); // @[FixedPointTypeClass.scala 21:58]
  assign _T_286 = $signed(io_in_bits_0) * $signed(io_weightMatrix_22_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_287 = $signed(io_in_bits_1) * $signed(io_weightMatrix_22_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_288 = $signed(io_in_bits_2) * $signed(io_weightMatrix_22_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_289 = $signed(io_in_bits_3) * $signed(io_weightMatrix_22_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_291 = $signed(_T_286) + $signed(_T_287); // @[FixedPointTypeClass.scala 21:58]
  assign _T_292 = $signed(_T_291); // @[FixedPointTypeClass.scala 21:58]
  assign _T_294 = $signed(_T_292) + $signed(_T_288); // @[FixedPointTypeClass.scala 21:58]
  assign _T_295 = $signed(_T_294); // @[FixedPointTypeClass.scala 21:58]
  assign _T_297 = $signed(_T_295) + $signed(_T_289); // @[FixedPointTypeClass.scala 21:58]
  assign _T_298 = $signed(_T_297); // @[FixedPointTypeClass.scala 21:58]
  assign _T_299 = $signed(io_in_bits_0) * $signed(io_weightMatrix_23_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_300 = $signed(io_in_bits_1) * $signed(io_weightMatrix_23_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_301 = $signed(io_in_bits_2) * $signed(io_weightMatrix_23_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_302 = $signed(io_in_bits_3) * $signed(io_weightMatrix_23_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_304 = $signed(_T_299) + $signed(_T_300); // @[FixedPointTypeClass.scala 21:58]
  assign _T_305 = $signed(_T_304); // @[FixedPointTypeClass.scala 21:58]
  assign _T_307 = $signed(_T_305) + $signed(_T_301); // @[FixedPointTypeClass.scala 21:58]
  assign _T_308 = $signed(_T_307); // @[FixedPointTypeClass.scala 21:58]
  assign _T_310 = $signed(_T_308) + $signed(_T_302); // @[FixedPointTypeClass.scala 21:58]
  assign _T_311 = $signed(_T_310); // @[FixedPointTypeClass.scala 21:58]
  assign _T_312 = $signed(io_in_bits_0) * $signed(io_weightMatrix_24_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_313 = $signed(io_in_bits_1) * $signed(io_weightMatrix_24_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_314 = $signed(io_in_bits_2) * $signed(io_weightMatrix_24_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_315 = $signed(io_in_bits_3) * $signed(io_weightMatrix_24_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_317 = $signed(_T_312) + $signed(_T_313); // @[FixedPointTypeClass.scala 21:58]
  assign _T_318 = $signed(_T_317); // @[FixedPointTypeClass.scala 21:58]
  assign _T_320 = $signed(_T_318) + $signed(_T_314); // @[FixedPointTypeClass.scala 21:58]
  assign _T_321 = $signed(_T_320); // @[FixedPointTypeClass.scala 21:58]
  assign _T_323 = $signed(_T_321) + $signed(_T_315); // @[FixedPointTypeClass.scala 21:58]
  assign _T_324 = $signed(_T_323); // @[FixedPointTypeClass.scala 21:58]
  assign _T_325 = $signed(io_in_bits_0) * $signed(io_weightMatrix_25_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_326 = $signed(io_in_bits_1) * $signed(io_weightMatrix_25_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_327 = $signed(io_in_bits_2) * $signed(io_weightMatrix_25_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_328 = $signed(io_in_bits_3) * $signed(io_weightMatrix_25_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_330 = $signed(_T_325) + $signed(_T_326); // @[FixedPointTypeClass.scala 21:58]
  assign _T_331 = $signed(_T_330); // @[FixedPointTypeClass.scala 21:58]
  assign _T_333 = $signed(_T_331) + $signed(_T_327); // @[FixedPointTypeClass.scala 21:58]
  assign _T_334 = $signed(_T_333); // @[FixedPointTypeClass.scala 21:58]
  assign _T_336 = $signed(_T_334) + $signed(_T_328); // @[FixedPointTypeClass.scala 21:58]
  assign _T_337 = $signed(_T_336); // @[FixedPointTypeClass.scala 21:58]
  assign _T_338 = $signed(io_in_bits_0) * $signed(io_weightMatrix_26_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_339 = $signed(io_in_bits_1) * $signed(io_weightMatrix_26_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_340 = $signed(io_in_bits_2) * $signed(io_weightMatrix_26_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_341 = $signed(io_in_bits_3) * $signed(io_weightMatrix_26_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_343 = $signed(_T_338) + $signed(_T_339); // @[FixedPointTypeClass.scala 21:58]
  assign _T_344 = $signed(_T_343); // @[FixedPointTypeClass.scala 21:58]
  assign _T_346 = $signed(_T_344) + $signed(_T_340); // @[FixedPointTypeClass.scala 21:58]
  assign _T_347 = $signed(_T_346); // @[FixedPointTypeClass.scala 21:58]
  assign _T_349 = $signed(_T_347) + $signed(_T_341); // @[FixedPointTypeClass.scala 21:58]
  assign _T_350 = $signed(_T_349); // @[FixedPointTypeClass.scala 21:58]
  assign _T_351 = $signed(io_in_bits_0) * $signed(io_weightMatrix_27_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_352 = $signed(io_in_bits_1) * $signed(io_weightMatrix_27_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_353 = $signed(io_in_bits_2) * $signed(io_weightMatrix_27_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_354 = $signed(io_in_bits_3) * $signed(io_weightMatrix_27_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_356 = $signed(_T_351) + $signed(_T_352); // @[FixedPointTypeClass.scala 21:58]
  assign _T_357 = $signed(_T_356); // @[FixedPointTypeClass.scala 21:58]
  assign _T_359 = $signed(_T_357) + $signed(_T_353); // @[FixedPointTypeClass.scala 21:58]
  assign _T_360 = $signed(_T_359); // @[FixedPointTypeClass.scala 21:58]
  assign _T_362 = $signed(_T_360) + $signed(_T_354); // @[FixedPointTypeClass.scala 21:58]
  assign _T_363 = $signed(_T_362); // @[FixedPointTypeClass.scala 21:58]
  assign _T_364 = $signed(io_in_bits_0) * $signed(io_weightMatrix_28_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_365 = $signed(io_in_bits_1) * $signed(io_weightMatrix_28_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_366 = $signed(io_in_bits_2) * $signed(io_weightMatrix_28_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_367 = $signed(io_in_bits_3) * $signed(io_weightMatrix_28_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_369 = $signed(_T_364) + $signed(_T_365); // @[FixedPointTypeClass.scala 21:58]
  assign _T_370 = $signed(_T_369); // @[FixedPointTypeClass.scala 21:58]
  assign _T_372 = $signed(_T_370) + $signed(_T_366); // @[FixedPointTypeClass.scala 21:58]
  assign _T_373 = $signed(_T_372); // @[FixedPointTypeClass.scala 21:58]
  assign _T_375 = $signed(_T_373) + $signed(_T_367); // @[FixedPointTypeClass.scala 21:58]
  assign _T_376 = $signed(_T_375); // @[FixedPointTypeClass.scala 21:58]
  assign _T_377 = $signed(io_in_bits_0) * $signed(io_weightMatrix_29_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_378 = $signed(io_in_bits_1) * $signed(io_weightMatrix_29_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_379 = $signed(io_in_bits_2) * $signed(io_weightMatrix_29_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_380 = $signed(io_in_bits_3) * $signed(io_weightMatrix_29_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_382 = $signed(_T_377) + $signed(_T_378); // @[FixedPointTypeClass.scala 21:58]
  assign _T_383 = $signed(_T_382); // @[FixedPointTypeClass.scala 21:58]
  assign _T_385 = $signed(_T_383) + $signed(_T_379); // @[FixedPointTypeClass.scala 21:58]
  assign _T_386 = $signed(_T_385); // @[FixedPointTypeClass.scala 21:58]
  assign _T_388 = $signed(_T_386) + $signed(_T_380); // @[FixedPointTypeClass.scala 21:58]
  assign _T_389 = $signed(_T_388); // @[FixedPointTypeClass.scala 21:58]
  assign _T_390 = $signed(io_in_bits_0) * $signed(io_weightMatrix_30_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_391 = $signed(io_in_bits_1) * $signed(io_weightMatrix_30_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_392 = $signed(io_in_bits_2) * $signed(io_weightMatrix_30_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_393 = $signed(io_in_bits_3) * $signed(io_weightMatrix_30_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_395 = $signed(_T_390) + $signed(_T_391); // @[FixedPointTypeClass.scala 21:58]
  assign _T_396 = $signed(_T_395); // @[FixedPointTypeClass.scala 21:58]
  assign _T_398 = $signed(_T_396) + $signed(_T_392); // @[FixedPointTypeClass.scala 21:58]
  assign _T_399 = $signed(_T_398); // @[FixedPointTypeClass.scala 21:58]
  assign _T_401 = $signed(_T_399) + $signed(_T_393); // @[FixedPointTypeClass.scala 21:58]
  assign _T_402 = $signed(_T_401); // @[FixedPointTypeClass.scala 21:58]
  assign _T_403 = $signed(io_in_bits_0) * $signed(io_weightMatrix_31_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_404 = $signed(io_in_bits_1) * $signed(io_weightMatrix_31_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_405 = $signed(io_in_bits_2) * $signed(io_weightMatrix_31_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_406 = $signed(io_in_bits_3) * $signed(io_weightMatrix_31_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_408 = $signed(_T_403) + $signed(_T_404); // @[FixedPointTypeClass.scala 21:58]
  assign _T_409 = $signed(_T_408); // @[FixedPointTypeClass.scala 21:58]
  assign _T_411 = $signed(_T_409) + $signed(_T_405); // @[FixedPointTypeClass.scala 21:58]
  assign _T_412 = $signed(_T_411); // @[FixedPointTypeClass.scala 21:58]
  assign _T_414 = $signed(_T_412) + $signed(_T_406); // @[FixedPointTypeClass.scala 21:58]
  assign _T_415 = $signed(_T_414); // @[FixedPointTypeClass.scala 21:58]
  assign _T_416 = $signed(io_in_bits_0) * $signed(io_weightMatrix_32_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_417 = $signed(io_in_bits_1) * $signed(io_weightMatrix_32_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_418 = $signed(io_in_bits_2) * $signed(io_weightMatrix_32_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_419 = $signed(io_in_bits_3) * $signed(io_weightMatrix_32_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_421 = $signed(_T_416) + $signed(_T_417); // @[FixedPointTypeClass.scala 21:58]
  assign _T_422 = $signed(_T_421); // @[FixedPointTypeClass.scala 21:58]
  assign _T_424 = $signed(_T_422) + $signed(_T_418); // @[FixedPointTypeClass.scala 21:58]
  assign _T_425 = $signed(_T_424); // @[FixedPointTypeClass.scala 21:58]
  assign _T_427 = $signed(_T_425) + $signed(_T_419); // @[FixedPointTypeClass.scala 21:58]
  assign _T_428 = $signed(_T_427); // @[FixedPointTypeClass.scala 21:58]
  assign _T_429 = $signed(io_in_bits_0) * $signed(io_weightMatrix_33_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_430 = $signed(io_in_bits_1) * $signed(io_weightMatrix_33_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_431 = $signed(io_in_bits_2) * $signed(io_weightMatrix_33_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_432 = $signed(io_in_bits_3) * $signed(io_weightMatrix_33_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_434 = $signed(_T_429) + $signed(_T_430); // @[FixedPointTypeClass.scala 21:58]
  assign _T_435 = $signed(_T_434); // @[FixedPointTypeClass.scala 21:58]
  assign _T_437 = $signed(_T_435) + $signed(_T_431); // @[FixedPointTypeClass.scala 21:58]
  assign _T_438 = $signed(_T_437); // @[FixedPointTypeClass.scala 21:58]
  assign _T_440 = $signed(_T_438) + $signed(_T_432); // @[FixedPointTypeClass.scala 21:58]
  assign _T_441 = $signed(_T_440); // @[FixedPointTypeClass.scala 21:58]
  assign _T_442 = $signed(io_in_bits_0) * $signed(io_weightMatrix_34_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_443 = $signed(io_in_bits_1) * $signed(io_weightMatrix_34_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_444 = $signed(io_in_bits_2) * $signed(io_weightMatrix_34_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_445 = $signed(io_in_bits_3) * $signed(io_weightMatrix_34_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_447 = $signed(_T_442) + $signed(_T_443); // @[FixedPointTypeClass.scala 21:58]
  assign _T_448 = $signed(_T_447); // @[FixedPointTypeClass.scala 21:58]
  assign _T_450 = $signed(_T_448) + $signed(_T_444); // @[FixedPointTypeClass.scala 21:58]
  assign _T_451 = $signed(_T_450); // @[FixedPointTypeClass.scala 21:58]
  assign _T_453 = $signed(_T_451) + $signed(_T_445); // @[FixedPointTypeClass.scala 21:58]
  assign _T_454 = $signed(_T_453); // @[FixedPointTypeClass.scala 21:58]
  assign _T_455 = $signed(io_in_bits_0) * $signed(io_weightMatrix_35_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_456 = $signed(io_in_bits_1) * $signed(io_weightMatrix_35_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_457 = $signed(io_in_bits_2) * $signed(io_weightMatrix_35_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_458 = $signed(io_in_bits_3) * $signed(io_weightMatrix_35_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_460 = $signed(_T_455) + $signed(_T_456); // @[FixedPointTypeClass.scala 21:58]
  assign _T_461 = $signed(_T_460); // @[FixedPointTypeClass.scala 21:58]
  assign _T_463 = $signed(_T_461) + $signed(_T_457); // @[FixedPointTypeClass.scala 21:58]
  assign _T_464 = $signed(_T_463); // @[FixedPointTypeClass.scala 21:58]
  assign _T_466 = $signed(_T_464) + $signed(_T_458); // @[FixedPointTypeClass.scala 21:58]
  assign _T_467 = $signed(_T_466); // @[FixedPointTypeClass.scala 21:58]
  assign _T_468 = $signed(io_in_bits_0) * $signed(io_weightMatrix_36_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_469 = $signed(io_in_bits_1) * $signed(io_weightMatrix_36_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_470 = $signed(io_in_bits_2) * $signed(io_weightMatrix_36_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_471 = $signed(io_in_bits_3) * $signed(io_weightMatrix_36_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_473 = $signed(_T_468) + $signed(_T_469); // @[FixedPointTypeClass.scala 21:58]
  assign _T_474 = $signed(_T_473); // @[FixedPointTypeClass.scala 21:58]
  assign _T_476 = $signed(_T_474) + $signed(_T_470); // @[FixedPointTypeClass.scala 21:58]
  assign _T_477 = $signed(_T_476); // @[FixedPointTypeClass.scala 21:58]
  assign _T_479 = $signed(_T_477) + $signed(_T_471); // @[FixedPointTypeClass.scala 21:58]
  assign _T_480 = $signed(_T_479); // @[FixedPointTypeClass.scala 21:58]
  assign _T_481 = $signed(io_in_bits_0) * $signed(io_weightMatrix_37_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_482 = $signed(io_in_bits_1) * $signed(io_weightMatrix_37_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_483 = $signed(io_in_bits_2) * $signed(io_weightMatrix_37_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_484 = $signed(io_in_bits_3) * $signed(io_weightMatrix_37_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_486 = $signed(_T_481) + $signed(_T_482); // @[FixedPointTypeClass.scala 21:58]
  assign _T_487 = $signed(_T_486); // @[FixedPointTypeClass.scala 21:58]
  assign _T_489 = $signed(_T_487) + $signed(_T_483); // @[FixedPointTypeClass.scala 21:58]
  assign _T_490 = $signed(_T_489); // @[FixedPointTypeClass.scala 21:58]
  assign _T_492 = $signed(_T_490) + $signed(_T_484); // @[FixedPointTypeClass.scala 21:58]
  assign _T_493 = $signed(_T_492); // @[FixedPointTypeClass.scala 21:58]
  assign _T_494 = $signed(io_in_bits_0) * $signed(io_weightMatrix_38_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_495 = $signed(io_in_bits_1) * $signed(io_weightMatrix_38_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_496 = $signed(io_in_bits_2) * $signed(io_weightMatrix_38_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_497 = $signed(io_in_bits_3) * $signed(io_weightMatrix_38_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_499 = $signed(_T_494) + $signed(_T_495); // @[FixedPointTypeClass.scala 21:58]
  assign _T_500 = $signed(_T_499); // @[FixedPointTypeClass.scala 21:58]
  assign _T_502 = $signed(_T_500) + $signed(_T_496); // @[FixedPointTypeClass.scala 21:58]
  assign _T_503 = $signed(_T_502); // @[FixedPointTypeClass.scala 21:58]
  assign _T_505 = $signed(_T_503) + $signed(_T_497); // @[FixedPointTypeClass.scala 21:58]
  assign _T_506 = $signed(_T_505); // @[FixedPointTypeClass.scala 21:58]
  assign _T_507 = $signed(io_in_bits_0) * $signed(io_weightMatrix_39_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_508 = $signed(io_in_bits_1) * $signed(io_weightMatrix_39_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_509 = $signed(io_in_bits_2) * $signed(io_weightMatrix_39_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_510 = $signed(io_in_bits_3) * $signed(io_weightMatrix_39_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_512 = $signed(_T_507) + $signed(_T_508); // @[FixedPointTypeClass.scala 21:58]
  assign _T_513 = $signed(_T_512); // @[FixedPointTypeClass.scala 21:58]
  assign _T_515 = $signed(_T_513) + $signed(_T_509); // @[FixedPointTypeClass.scala 21:58]
  assign _T_516 = $signed(_T_515); // @[FixedPointTypeClass.scala 21:58]
  assign _T_518 = $signed(_T_516) + $signed(_T_510); // @[FixedPointTypeClass.scala 21:58]
  assign _T_519 = $signed(_T_518); // @[FixedPointTypeClass.scala 21:58]
  assign _T_520 = $signed(io_in_bits_0) * $signed(io_weightMatrix_40_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_521 = $signed(io_in_bits_1) * $signed(io_weightMatrix_40_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_522 = $signed(io_in_bits_2) * $signed(io_weightMatrix_40_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_523 = $signed(io_in_bits_3) * $signed(io_weightMatrix_40_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_525 = $signed(_T_520) + $signed(_T_521); // @[FixedPointTypeClass.scala 21:58]
  assign _T_526 = $signed(_T_525); // @[FixedPointTypeClass.scala 21:58]
  assign _T_528 = $signed(_T_526) + $signed(_T_522); // @[FixedPointTypeClass.scala 21:58]
  assign _T_529 = $signed(_T_528); // @[FixedPointTypeClass.scala 21:58]
  assign _T_531 = $signed(_T_529) + $signed(_T_523); // @[FixedPointTypeClass.scala 21:58]
  assign _T_532 = $signed(_T_531); // @[FixedPointTypeClass.scala 21:58]
  assign _T_533 = $signed(io_in_bits_0) * $signed(io_weightMatrix_41_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_534 = $signed(io_in_bits_1) * $signed(io_weightMatrix_41_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_535 = $signed(io_in_bits_2) * $signed(io_weightMatrix_41_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_536 = $signed(io_in_bits_3) * $signed(io_weightMatrix_41_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_538 = $signed(_T_533) + $signed(_T_534); // @[FixedPointTypeClass.scala 21:58]
  assign _T_539 = $signed(_T_538); // @[FixedPointTypeClass.scala 21:58]
  assign _T_541 = $signed(_T_539) + $signed(_T_535); // @[FixedPointTypeClass.scala 21:58]
  assign _T_542 = $signed(_T_541); // @[FixedPointTypeClass.scala 21:58]
  assign _T_544 = $signed(_T_542) + $signed(_T_536); // @[FixedPointTypeClass.scala 21:58]
  assign _T_545 = $signed(_T_544); // @[FixedPointTypeClass.scala 21:58]
  assign _T_546 = $signed(io_in_bits_0) * $signed(io_weightMatrix_42_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_547 = $signed(io_in_bits_1) * $signed(io_weightMatrix_42_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_548 = $signed(io_in_bits_2) * $signed(io_weightMatrix_42_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_549 = $signed(io_in_bits_3) * $signed(io_weightMatrix_42_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_551 = $signed(_T_546) + $signed(_T_547); // @[FixedPointTypeClass.scala 21:58]
  assign _T_552 = $signed(_T_551); // @[FixedPointTypeClass.scala 21:58]
  assign _T_554 = $signed(_T_552) + $signed(_T_548); // @[FixedPointTypeClass.scala 21:58]
  assign _T_555 = $signed(_T_554); // @[FixedPointTypeClass.scala 21:58]
  assign _T_557 = $signed(_T_555) + $signed(_T_549); // @[FixedPointTypeClass.scala 21:58]
  assign _T_558 = $signed(_T_557); // @[FixedPointTypeClass.scala 21:58]
  assign _T_559 = $signed(io_in_bits_0) * $signed(io_weightMatrix_43_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_560 = $signed(io_in_bits_1) * $signed(io_weightMatrix_43_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_561 = $signed(io_in_bits_2) * $signed(io_weightMatrix_43_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_562 = $signed(io_in_bits_3) * $signed(io_weightMatrix_43_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_564 = $signed(_T_559) + $signed(_T_560); // @[FixedPointTypeClass.scala 21:58]
  assign _T_565 = $signed(_T_564); // @[FixedPointTypeClass.scala 21:58]
  assign _T_567 = $signed(_T_565) + $signed(_T_561); // @[FixedPointTypeClass.scala 21:58]
  assign _T_568 = $signed(_T_567); // @[FixedPointTypeClass.scala 21:58]
  assign _T_570 = $signed(_T_568) + $signed(_T_562); // @[FixedPointTypeClass.scala 21:58]
  assign _T_571 = $signed(_T_570); // @[FixedPointTypeClass.scala 21:58]
  assign _T_572 = $signed(io_in_bits_0) * $signed(io_weightMatrix_44_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_573 = $signed(io_in_bits_1) * $signed(io_weightMatrix_44_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_574 = $signed(io_in_bits_2) * $signed(io_weightMatrix_44_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_575 = $signed(io_in_bits_3) * $signed(io_weightMatrix_44_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_577 = $signed(_T_572) + $signed(_T_573); // @[FixedPointTypeClass.scala 21:58]
  assign _T_578 = $signed(_T_577); // @[FixedPointTypeClass.scala 21:58]
  assign _T_580 = $signed(_T_578) + $signed(_T_574); // @[FixedPointTypeClass.scala 21:58]
  assign _T_581 = $signed(_T_580); // @[FixedPointTypeClass.scala 21:58]
  assign _T_583 = $signed(_T_581) + $signed(_T_575); // @[FixedPointTypeClass.scala 21:58]
  assign _T_584 = $signed(_T_583); // @[FixedPointTypeClass.scala 21:58]
  assign _T_585 = $signed(io_in_bits_0) * $signed(io_weightMatrix_45_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_586 = $signed(io_in_bits_1) * $signed(io_weightMatrix_45_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_587 = $signed(io_in_bits_2) * $signed(io_weightMatrix_45_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_588 = $signed(io_in_bits_3) * $signed(io_weightMatrix_45_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_590 = $signed(_T_585) + $signed(_T_586); // @[FixedPointTypeClass.scala 21:58]
  assign _T_591 = $signed(_T_590); // @[FixedPointTypeClass.scala 21:58]
  assign _T_593 = $signed(_T_591) + $signed(_T_587); // @[FixedPointTypeClass.scala 21:58]
  assign _T_594 = $signed(_T_593); // @[FixedPointTypeClass.scala 21:58]
  assign _T_596 = $signed(_T_594) + $signed(_T_588); // @[FixedPointTypeClass.scala 21:58]
  assign _T_597 = $signed(_T_596); // @[FixedPointTypeClass.scala 21:58]
  assign _T_598 = $signed(io_in_bits_0) * $signed(io_weightMatrix_46_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_599 = $signed(io_in_bits_1) * $signed(io_weightMatrix_46_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_600 = $signed(io_in_bits_2) * $signed(io_weightMatrix_46_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_601 = $signed(io_in_bits_3) * $signed(io_weightMatrix_46_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_603 = $signed(_T_598) + $signed(_T_599); // @[FixedPointTypeClass.scala 21:58]
  assign _T_604 = $signed(_T_603); // @[FixedPointTypeClass.scala 21:58]
  assign _T_606 = $signed(_T_604) + $signed(_T_600); // @[FixedPointTypeClass.scala 21:58]
  assign _T_607 = $signed(_T_606); // @[FixedPointTypeClass.scala 21:58]
  assign _T_609 = $signed(_T_607) + $signed(_T_601); // @[FixedPointTypeClass.scala 21:58]
  assign _T_610 = $signed(_T_609); // @[FixedPointTypeClass.scala 21:58]
  assign _T_611 = $signed(io_in_bits_0) * $signed(io_weightMatrix_47_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_612 = $signed(io_in_bits_1) * $signed(io_weightMatrix_47_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_613 = $signed(io_in_bits_2) * $signed(io_weightMatrix_47_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_614 = $signed(io_in_bits_3) * $signed(io_weightMatrix_47_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_616 = $signed(_T_611) + $signed(_T_612); // @[FixedPointTypeClass.scala 21:58]
  assign _T_617 = $signed(_T_616); // @[FixedPointTypeClass.scala 21:58]
  assign _T_619 = $signed(_T_617) + $signed(_T_613); // @[FixedPointTypeClass.scala 21:58]
  assign _T_620 = $signed(_T_619); // @[FixedPointTypeClass.scala 21:58]
  assign _T_622 = $signed(_T_620) + $signed(_T_614); // @[FixedPointTypeClass.scala 21:58]
  assign _T_623 = $signed(_T_622); // @[FixedPointTypeClass.scala 21:58]
  assign _T_624 = $signed(io_in_bits_0) * $signed(io_weightMatrix_48_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_625 = $signed(io_in_bits_1) * $signed(io_weightMatrix_48_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_626 = $signed(io_in_bits_2) * $signed(io_weightMatrix_48_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_627 = $signed(io_in_bits_3) * $signed(io_weightMatrix_48_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_629 = $signed(_T_624) + $signed(_T_625); // @[FixedPointTypeClass.scala 21:58]
  assign _T_630 = $signed(_T_629); // @[FixedPointTypeClass.scala 21:58]
  assign _T_632 = $signed(_T_630) + $signed(_T_626); // @[FixedPointTypeClass.scala 21:58]
  assign _T_633 = $signed(_T_632); // @[FixedPointTypeClass.scala 21:58]
  assign _T_635 = $signed(_T_633) + $signed(_T_627); // @[FixedPointTypeClass.scala 21:58]
  assign _T_636 = $signed(_T_635); // @[FixedPointTypeClass.scala 21:58]
  assign _T_637 = $signed(io_in_bits_0) * $signed(io_weightMatrix_49_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_638 = $signed(io_in_bits_1) * $signed(io_weightMatrix_49_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_639 = $signed(io_in_bits_2) * $signed(io_weightMatrix_49_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_640 = $signed(io_in_bits_3) * $signed(io_weightMatrix_49_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_642 = $signed(_T_637) + $signed(_T_638); // @[FixedPointTypeClass.scala 21:58]
  assign _T_643 = $signed(_T_642); // @[FixedPointTypeClass.scala 21:58]
  assign _T_645 = $signed(_T_643) + $signed(_T_639); // @[FixedPointTypeClass.scala 21:58]
  assign _T_646 = $signed(_T_645); // @[FixedPointTypeClass.scala 21:58]
  assign _T_648 = $signed(_T_646) + $signed(_T_640); // @[FixedPointTypeClass.scala 21:58]
  assign _T_649 = $signed(_T_648); // @[FixedPointTypeClass.scala 21:58]
  assign _T_650 = $signed(io_in_bits_0) * $signed(io_weightMatrix_50_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_651 = $signed(io_in_bits_1) * $signed(io_weightMatrix_50_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_652 = $signed(io_in_bits_2) * $signed(io_weightMatrix_50_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_653 = $signed(io_in_bits_3) * $signed(io_weightMatrix_50_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_655 = $signed(_T_650) + $signed(_T_651); // @[FixedPointTypeClass.scala 21:58]
  assign _T_656 = $signed(_T_655); // @[FixedPointTypeClass.scala 21:58]
  assign _T_658 = $signed(_T_656) + $signed(_T_652); // @[FixedPointTypeClass.scala 21:58]
  assign _T_659 = $signed(_T_658); // @[FixedPointTypeClass.scala 21:58]
  assign _T_661 = $signed(_T_659) + $signed(_T_653); // @[FixedPointTypeClass.scala 21:58]
  assign _T_662 = $signed(_T_661); // @[FixedPointTypeClass.scala 21:58]
  assign _T_663 = $signed(io_in_bits_0) * $signed(io_weightMatrix_51_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_664 = $signed(io_in_bits_1) * $signed(io_weightMatrix_51_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_665 = $signed(io_in_bits_2) * $signed(io_weightMatrix_51_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_666 = $signed(io_in_bits_3) * $signed(io_weightMatrix_51_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_668 = $signed(_T_663) + $signed(_T_664); // @[FixedPointTypeClass.scala 21:58]
  assign _T_669 = $signed(_T_668); // @[FixedPointTypeClass.scala 21:58]
  assign _T_671 = $signed(_T_669) + $signed(_T_665); // @[FixedPointTypeClass.scala 21:58]
  assign _T_672 = $signed(_T_671); // @[FixedPointTypeClass.scala 21:58]
  assign _T_674 = $signed(_T_672) + $signed(_T_666); // @[FixedPointTypeClass.scala 21:58]
  assign _T_675 = $signed(_T_674); // @[FixedPointTypeClass.scala 21:58]
  assign _T_676 = $signed(io_in_bits_0) * $signed(io_weightMatrix_52_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_677 = $signed(io_in_bits_1) * $signed(io_weightMatrix_52_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_678 = $signed(io_in_bits_2) * $signed(io_weightMatrix_52_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_679 = $signed(io_in_bits_3) * $signed(io_weightMatrix_52_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_681 = $signed(_T_676) + $signed(_T_677); // @[FixedPointTypeClass.scala 21:58]
  assign _T_682 = $signed(_T_681); // @[FixedPointTypeClass.scala 21:58]
  assign _T_684 = $signed(_T_682) + $signed(_T_678); // @[FixedPointTypeClass.scala 21:58]
  assign _T_685 = $signed(_T_684); // @[FixedPointTypeClass.scala 21:58]
  assign _T_687 = $signed(_T_685) + $signed(_T_679); // @[FixedPointTypeClass.scala 21:58]
  assign _T_688 = $signed(_T_687); // @[FixedPointTypeClass.scala 21:58]
  assign _T_689 = $signed(io_in_bits_0) * $signed(io_weightMatrix_53_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_690 = $signed(io_in_bits_1) * $signed(io_weightMatrix_53_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_691 = $signed(io_in_bits_2) * $signed(io_weightMatrix_53_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_692 = $signed(io_in_bits_3) * $signed(io_weightMatrix_53_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_694 = $signed(_T_689) + $signed(_T_690); // @[FixedPointTypeClass.scala 21:58]
  assign _T_695 = $signed(_T_694); // @[FixedPointTypeClass.scala 21:58]
  assign _T_697 = $signed(_T_695) + $signed(_T_691); // @[FixedPointTypeClass.scala 21:58]
  assign _T_698 = $signed(_T_697); // @[FixedPointTypeClass.scala 21:58]
  assign _T_700 = $signed(_T_698) + $signed(_T_692); // @[FixedPointTypeClass.scala 21:58]
  assign _T_701 = $signed(_T_700); // @[FixedPointTypeClass.scala 21:58]
  assign _T_702 = $signed(io_in_bits_0) * $signed(io_weightMatrix_54_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_703 = $signed(io_in_bits_1) * $signed(io_weightMatrix_54_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_704 = $signed(io_in_bits_2) * $signed(io_weightMatrix_54_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_705 = $signed(io_in_bits_3) * $signed(io_weightMatrix_54_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_707 = $signed(_T_702) + $signed(_T_703); // @[FixedPointTypeClass.scala 21:58]
  assign _T_708 = $signed(_T_707); // @[FixedPointTypeClass.scala 21:58]
  assign _T_710 = $signed(_T_708) + $signed(_T_704); // @[FixedPointTypeClass.scala 21:58]
  assign _T_711 = $signed(_T_710); // @[FixedPointTypeClass.scala 21:58]
  assign _T_713 = $signed(_T_711) + $signed(_T_705); // @[FixedPointTypeClass.scala 21:58]
  assign _T_714 = $signed(_T_713); // @[FixedPointTypeClass.scala 21:58]
  assign _T_715 = $signed(io_in_bits_0) * $signed(io_weightMatrix_55_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_716 = $signed(io_in_bits_1) * $signed(io_weightMatrix_55_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_717 = $signed(io_in_bits_2) * $signed(io_weightMatrix_55_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_718 = $signed(io_in_bits_3) * $signed(io_weightMatrix_55_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_720 = $signed(_T_715) + $signed(_T_716); // @[FixedPointTypeClass.scala 21:58]
  assign _T_721 = $signed(_T_720); // @[FixedPointTypeClass.scala 21:58]
  assign _T_723 = $signed(_T_721) + $signed(_T_717); // @[FixedPointTypeClass.scala 21:58]
  assign _T_724 = $signed(_T_723); // @[FixedPointTypeClass.scala 21:58]
  assign _T_726 = $signed(_T_724) + $signed(_T_718); // @[FixedPointTypeClass.scala 21:58]
  assign _T_727 = $signed(_T_726); // @[FixedPointTypeClass.scala 21:58]
  assign _T_728 = $signed(io_in_bits_0) * $signed(io_weightMatrix_56_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_729 = $signed(io_in_bits_1) * $signed(io_weightMatrix_56_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_730 = $signed(io_in_bits_2) * $signed(io_weightMatrix_56_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_731 = $signed(io_in_bits_3) * $signed(io_weightMatrix_56_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_733 = $signed(_T_728) + $signed(_T_729); // @[FixedPointTypeClass.scala 21:58]
  assign _T_734 = $signed(_T_733); // @[FixedPointTypeClass.scala 21:58]
  assign _T_736 = $signed(_T_734) + $signed(_T_730); // @[FixedPointTypeClass.scala 21:58]
  assign _T_737 = $signed(_T_736); // @[FixedPointTypeClass.scala 21:58]
  assign _T_739 = $signed(_T_737) + $signed(_T_731); // @[FixedPointTypeClass.scala 21:58]
  assign _T_740 = $signed(_T_739); // @[FixedPointTypeClass.scala 21:58]
  assign _T_741 = $signed(io_in_bits_0) * $signed(io_weightMatrix_57_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_742 = $signed(io_in_bits_1) * $signed(io_weightMatrix_57_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_743 = $signed(io_in_bits_2) * $signed(io_weightMatrix_57_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_744 = $signed(io_in_bits_3) * $signed(io_weightMatrix_57_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_746 = $signed(_T_741) + $signed(_T_742); // @[FixedPointTypeClass.scala 21:58]
  assign _T_747 = $signed(_T_746); // @[FixedPointTypeClass.scala 21:58]
  assign _T_749 = $signed(_T_747) + $signed(_T_743); // @[FixedPointTypeClass.scala 21:58]
  assign _T_750 = $signed(_T_749); // @[FixedPointTypeClass.scala 21:58]
  assign _T_752 = $signed(_T_750) + $signed(_T_744); // @[FixedPointTypeClass.scala 21:58]
  assign _T_753 = $signed(_T_752); // @[FixedPointTypeClass.scala 21:58]
  assign _T_754 = $signed(io_in_bits_0) * $signed(io_weightMatrix_58_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_755 = $signed(io_in_bits_1) * $signed(io_weightMatrix_58_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_756 = $signed(io_in_bits_2) * $signed(io_weightMatrix_58_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_757 = $signed(io_in_bits_3) * $signed(io_weightMatrix_58_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_759 = $signed(_T_754) + $signed(_T_755); // @[FixedPointTypeClass.scala 21:58]
  assign _T_760 = $signed(_T_759); // @[FixedPointTypeClass.scala 21:58]
  assign _T_762 = $signed(_T_760) + $signed(_T_756); // @[FixedPointTypeClass.scala 21:58]
  assign _T_763 = $signed(_T_762); // @[FixedPointTypeClass.scala 21:58]
  assign _T_765 = $signed(_T_763) + $signed(_T_757); // @[FixedPointTypeClass.scala 21:58]
  assign _T_766 = $signed(_T_765); // @[FixedPointTypeClass.scala 21:58]
  assign _T_767 = $signed(io_in_bits_0) * $signed(io_weightMatrix_59_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_768 = $signed(io_in_bits_1) * $signed(io_weightMatrix_59_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_769 = $signed(io_in_bits_2) * $signed(io_weightMatrix_59_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_770 = $signed(io_in_bits_3) * $signed(io_weightMatrix_59_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_772 = $signed(_T_767) + $signed(_T_768); // @[FixedPointTypeClass.scala 21:58]
  assign _T_773 = $signed(_T_772); // @[FixedPointTypeClass.scala 21:58]
  assign _T_775 = $signed(_T_773) + $signed(_T_769); // @[FixedPointTypeClass.scala 21:58]
  assign _T_776 = $signed(_T_775); // @[FixedPointTypeClass.scala 21:58]
  assign _T_778 = $signed(_T_776) + $signed(_T_770); // @[FixedPointTypeClass.scala 21:58]
  assign _T_779 = $signed(_T_778); // @[FixedPointTypeClass.scala 21:58]
  assign _T_780 = $signed(io_in_bits_0) * $signed(io_weightMatrix_60_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_781 = $signed(io_in_bits_1) * $signed(io_weightMatrix_60_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_782 = $signed(io_in_bits_2) * $signed(io_weightMatrix_60_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_783 = $signed(io_in_bits_3) * $signed(io_weightMatrix_60_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_785 = $signed(_T_780) + $signed(_T_781); // @[FixedPointTypeClass.scala 21:58]
  assign _T_786 = $signed(_T_785); // @[FixedPointTypeClass.scala 21:58]
  assign _T_788 = $signed(_T_786) + $signed(_T_782); // @[FixedPointTypeClass.scala 21:58]
  assign _T_789 = $signed(_T_788); // @[FixedPointTypeClass.scala 21:58]
  assign _T_791 = $signed(_T_789) + $signed(_T_783); // @[FixedPointTypeClass.scala 21:58]
  assign _T_792 = $signed(_T_791); // @[FixedPointTypeClass.scala 21:58]
  assign _T_793 = $signed(io_in_bits_0) * $signed(io_weightMatrix_61_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_794 = $signed(io_in_bits_1) * $signed(io_weightMatrix_61_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_795 = $signed(io_in_bits_2) * $signed(io_weightMatrix_61_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_796 = $signed(io_in_bits_3) * $signed(io_weightMatrix_61_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_798 = $signed(_T_793) + $signed(_T_794); // @[FixedPointTypeClass.scala 21:58]
  assign _T_799 = $signed(_T_798); // @[FixedPointTypeClass.scala 21:58]
  assign _T_801 = $signed(_T_799) + $signed(_T_795); // @[FixedPointTypeClass.scala 21:58]
  assign _T_802 = $signed(_T_801); // @[FixedPointTypeClass.scala 21:58]
  assign _T_804 = $signed(_T_802) + $signed(_T_796); // @[FixedPointTypeClass.scala 21:58]
  assign _T_805 = $signed(_T_804); // @[FixedPointTypeClass.scala 21:58]
  assign _T_806 = $signed(io_in_bits_0) * $signed(io_weightMatrix_62_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_807 = $signed(io_in_bits_1) * $signed(io_weightMatrix_62_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_808 = $signed(io_in_bits_2) * $signed(io_weightMatrix_62_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_809 = $signed(io_in_bits_3) * $signed(io_weightMatrix_62_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_811 = $signed(_T_806) + $signed(_T_807); // @[FixedPointTypeClass.scala 21:58]
  assign _T_812 = $signed(_T_811); // @[FixedPointTypeClass.scala 21:58]
  assign _T_814 = $signed(_T_812) + $signed(_T_808); // @[FixedPointTypeClass.scala 21:58]
  assign _T_815 = $signed(_T_814); // @[FixedPointTypeClass.scala 21:58]
  assign _T_817 = $signed(_T_815) + $signed(_T_809); // @[FixedPointTypeClass.scala 21:58]
  assign _T_818 = $signed(_T_817); // @[FixedPointTypeClass.scala 21:58]
  assign _T_819 = $signed(io_in_bits_0) * $signed(io_weightMatrix_63_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_820 = $signed(io_in_bits_1) * $signed(io_weightMatrix_63_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_821 = $signed(io_in_bits_2) * $signed(io_weightMatrix_63_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_822 = $signed(io_in_bits_3) * $signed(io_weightMatrix_63_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_824 = $signed(_T_819) + $signed(_T_820); // @[FixedPointTypeClass.scala 21:58]
  assign _T_825 = $signed(_T_824); // @[FixedPointTypeClass.scala 21:58]
  assign _T_827 = $signed(_T_825) + $signed(_T_821); // @[FixedPointTypeClass.scala 21:58]
  assign _T_828 = $signed(_T_827); // @[FixedPointTypeClass.scala 21:58]
  assign _T_830 = $signed(_T_828) + $signed(_T_822); // @[FixedPointTypeClass.scala 21:58]
  assign _T_831 = $signed(_T_830); // @[FixedPointTypeClass.scala 21:58]
  assign _T_832 = $signed(io_in_bits_0) * $signed(io_weightMatrix_64_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_833 = $signed(io_in_bits_1) * $signed(io_weightMatrix_64_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_834 = $signed(io_in_bits_2) * $signed(io_weightMatrix_64_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_835 = $signed(io_in_bits_3) * $signed(io_weightMatrix_64_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_837 = $signed(_T_832) + $signed(_T_833); // @[FixedPointTypeClass.scala 21:58]
  assign _T_838 = $signed(_T_837); // @[FixedPointTypeClass.scala 21:58]
  assign _T_840 = $signed(_T_838) + $signed(_T_834); // @[FixedPointTypeClass.scala 21:58]
  assign _T_841 = $signed(_T_840); // @[FixedPointTypeClass.scala 21:58]
  assign _T_843 = $signed(_T_841) + $signed(_T_835); // @[FixedPointTypeClass.scala 21:58]
  assign _T_844 = $signed(_T_843); // @[FixedPointTypeClass.scala 21:58]
  assign _T_845 = $signed(io_in_bits_0) * $signed(io_weightMatrix_65_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_846 = $signed(io_in_bits_1) * $signed(io_weightMatrix_65_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_847 = $signed(io_in_bits_2) * $signed(io_weightMatrix_65_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_848 = $signed(io_in_bits_3) * $signed(io_weightMatrix_65_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_850 = $signed(_T_845) + $signed(_T_846); // @[FixedPointTypeClass.scala 21:58]
  assign _T_851 = $signed(_T_850); // @[FixedPointTypeClass.scala 21:58]
  assign _T_853 = $signed(_T_851) + $signed(_T_847); // @[FixedPointTypeClass.scala 21:58]
  assign _T_854 = $signed(_T_853); // @[FixedPointTypeClass.scala 21:58]
  assign _T_856 = $signed(_T_854) + $signed(_T_848); // @[FixedPointTypeClass.scala 21:58]
  assign _T_857 = $signed(_T_856); // @[FixedPointTypeClass.scala 21:58]
  assign _T_858 = $signed(io_in_bits_0) * $signed(io_weightMatrix_66_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_859 = $signed(io_in_bits_1) * $signed(io_weightMatrix_66_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_860 = $signed(io_in_bits_2) * $signed(io_weightMatrix_66_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_861 = $signed(io_in_bits_3) * $signed(io_weightMatrix_66_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_863 = $signed(_T_858) + $signed(_T_859); // @[FixedPointTypeClass.scala 21:58]
  assign _T_864 = $signed(_T_863); // @[FixedPointTypeClass.scala 21:58]
  assign _T_866 = $signed(_T_864) + $signed(_T_860); // @[FixedPointTypeClass.scala 21:58]
  assign _T_867 = $signed(_T_866); // @[FixedPointTypeClass.scala 21:58]
  assign _T_869 = $signed(_T_867) + $signed(_T_861); // @[FixedPointTypeClass.scala 21:58]
  assign _T_870 = $signed(_T_869); // @[FixedPointTypeClass.scala 21:58]
  assign _T_871 = $signed(io_in_bits_0) * $signed(io_weightMatrix_67_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_872 = $signed(io_in_bits_1) * $signed(io_weightMatrix_67_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_873 = $signed(io_in_bits_2) * $signed(io_weightMatrix_67_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_874 = $signed(io_in_bits_3) * $signed(io_weightMatrix_67_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_876 = $signed(_T_871) + $signed(_T_872); // @[FixedPointTypeClass.scala 21:58]
  assign _T_877 = $signed(_T_876); // @[FixedPointTypeClass.scala 21:58]
  assign _T_879 = $signed(_T_877) + $signed(_T_873); // @[FixedPointTypeClass.scala 21:58]
  assign _T_880 = $signed(_T_879); // @[FixedPointTypeClass.scala 21:58]
  assign _T_882 = $signed(_T_880) + $signed(_T_874); // @[FixedPointTypeClass.scala 21:58]
  assign _T_883 = $signed(_T_882); // @[FixedPointTypeClass.scala 21:58]
  assign _T_884 = $signed(io_in_bits_0) * $signed(io_weightMatrix_68_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_885 = $signed(io_in_bits_1) * $signed(io_weightMatrix_68_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_886 = $signed(io_in_bits_2) * $signed(io_weightMatrix_68_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_887 = $signed(io_in_bits_3) * $signed(io_weightMatrix_68_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_889 = $signed(_T_884) + $signed(_T_885); // @[FixedPointTypeClass.scala 21:58]
  assign _T_890 = $signed(_T_889); // @[FixedPointTypeClass.scala 21:58]
  assign _T_892 = $signed(_T_890) + $signed(_T_886); // @[FixedPointTypeClass.scala 21:58]
  assign _T_893 = $signed(_T_892); // @[FixedPointTypeClass.scala 21:58]
  assign _T_895 = $signed(_T_893) + $signed(_T_887); // @[FixedPointTypeClass.scala 21:58]
  assign _T_896 = $signed(_T_895); // @[FixedPointTypeClass.scala 21:58]
  assign _T_897 = $signed(io_in_bits_0) * $signed(io_weightMatrix_69_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_898 = $signed(io_in_bits_1) * $signed(io_weightMatrix_69_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_899 = $signed(io_in_bits_2) * $signed(io_weightMatrix_69_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_900 = $signed(io_in_bits_3) * $signed(io_weightMatrix_69_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_902 = $signed(_T_897) + $signed(_T_898); // @[FixedPointTypeClass.scala 21:58]
  assign _T_903 = $signed(_T_902); // @[FixedPointTypeClass.scala 21:58]
  assign _T_905 = $signed(_T_903) + $signed(_T_899); // @[FixedPointTypeClass.scala 21:58]
  assign _T_906 = $signed(_T_905); // @[FixedPointTypeClass.scala 21:58]
  assign _T_908 = $signed(_T_906) + $signed(_T_900); // @[FixedPointTypeClass.scala 21:58]
  assign _T_909 = $signed(_T_908); // @[FixedPointTypeClass.scala 21:58]
  assign _T_910 = $signed(io_in_bits_0) * $signed(io_weightMatrix_70_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_911 = $signed(io_in_bits_1) * $signed(io_weightMatrix_70_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_912 = $signed(io_in_bits_2) * $signed(io_weightMatrix_70_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_913 = $signed(io_in_bits_3) * $signed(io_weightMatrix_70_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_915 = $signed(_T_910) + $signed(_T_911); // @[FixedPointTypeClass.scala 21:58]
  assign _T_916 = $signed(_T_915); // @[FixedPointTypeClass.scala 21:58]
  assign _T_918 = $signed(_T_916) + $signed(_T_912); // @[FixedPointTypeClass.scala 21:58]
  assign _T_919 = $signed(_T_918); // @[FixedPointTypeClass.scala 21:58]
  assign _T_921 = $signed(_T_919) + $signed(_T_913); // @[FixedPointTypeClass.scala 21:58]
  assign _T_922 = $signed(_T_921); // @[FixedPointTypeClass.scala 21:58]
  assign _T_923 = $signed(io_in_bits_0) * $signed(io_weightMatrix_71_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_924 = $signed(io_in_bits_1) * $signed(io_weightMatrix_71_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_925 = $signed(io_in_bits_2) * $signed(io_weightMatrix_71_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_926 = $signed(io_in_bits_3) * $signed(io_weightMatrix_71_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_928 = $signed(_T_923) + $signed(_T_924); // @[FixedPointTypeClass.scala 21:58]
  assign _T_929 = $signed(_T_928); // @[FixedPointTypeClass.scala 21:58]
  assign _T_931 = $signed(_T_929) + $signed(_T_925); // @[FixedPointTypeClass.scala 21:58]
  assign _T_932 = $signed(_T_931); // @[FixedPointTypeClass.scala 21:58]
  assign _T_934 = $signed(_T_932) + $signed(_T_926); // @[FixedPointTypeClass.scala 21:58]
  assign _T_935 = $signed(_T_934); // @[FixedPointTypeClass.scala 21:58]
  assign _T_936 = $signed(io_in_bits_0) * $signed(io_weightMatrix_72_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_937 = $signed(io_in_bits_1) * $signed(io_weightMatrix_72_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_938 = $signed(io_in_bits_2) * $signed(io_weightMatrix_72_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_939 = $signed(io_in_bits_3) * $signed(io_weightMatrix_72_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_941 = $signed(_T_936) + $signed(_T_937); // @[FixedPointTypeClass.scala 21:58]
  assign _T_942 = $signed(_T_941); // @[FixedPointTypeClass.scala 21:58]
  assign _T_944 = $signed(_T_942) + $signed(_T_938); // @[FixedPointTypeClass.scala 21:58]
  assign _T_945 = $signed(_T_944); // @[FixedPointTypeClass.scala 21:58]
  assign _T_947 = $signed(_T_945) + $signed(_T_939); // @[FixedPointTypeClass.scala 21:58]
  assign _T_948 = $signed(_T_947); // @[FixedPointTypeClass.scala 21:58]
  assign _T_949 = $signed(io_in_bits_0) * $signed(io_weightMatrix_73_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_950 = $signed(io_in_bits_1) * $signed(io_weightMatrix_73_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_951 = $signed(io_in_bits_2) * $signed(io_weightMatrix_73_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_952 = $signed(io_in_bits_3) * $signed(io_weightMatrix_73_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_954 = $signed(_T_949) + $signed(_T_950); // @[FixedPointTypeClass.scala 21:58]
  assign _T_955 = $signed(_T_954); // @[FixedPointTypeClass.scala 21:58]
  assign _T_957 = $signed(_T_955) + $signed(_T_951); // @[FixedPointTypeClass.scala 21:58]
  assign _T_958 = $signed(_T_957); // @[FixedPointTypeClass.scala 21:58]
  assign _T_960 = $signed(_T_958) + $signed(_T_952); // @[FixedPointTypeClass.scala 21:58]
  assign _T_961 = $signed(_T_960); // @[FixedPointTypeClass.scala 21:58]
  assign _T_962 = $signed(io_in_bits_0) * $signed(io_weightMatrix_74_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_963 = $signed(io_in_bits_1) * $signed(io_weightMatrix_74_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_964 = $signed(io_in_bits_2) * $signed(io_weightMatrix_74_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_965 = $signed(io_in_bits_3) * $signed(io_weightMatrix_74_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_967 = $signed(_T_962) + $signed(_T_963); // @[FixedPointTypeClass.scala 21:58]
  assign _T_968 = $signed(_T_967); // @[FixedPointTypeClass.scala 21:58]
  assign _T_970 = $signed(_T_968) + $signed(_T_964); // @[FixedPointTypeClass.scala 21:58]
  assign _T_971 = $signed(_T_970); // @[FixedPointTypeClass.scala 21:58]
  assign _T_973 = $signed(_T_971) + $signed(_T_965); // @[FixedPointTypeClass.scala 21:58]
  assign _T_974 = $signed(_T_973); // @[FixedPointTypeClass.scala 21:58]
  assign _T_975 = $signed(io_in_bits_0) * $signed(io_weightMatrix_75_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_976 = $signed(io_in_bits_1) * $signed(io_weightMatrix_75_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_977 = $signed(io_in_bits_2) * $signed(io_weightMatrix_75_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_978 = $signed(io_in_bits_3) * $signed(io_weightMatrix_75_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_980 = $signed(_T_975) + $signed(_T_976); // @[FixedPointTypeClass.scala 21:58]
  assign _T_981 = $signed(_T_980); // @[FixedPointTypeClass.scala 21:58]
  assign _T_983 = $signed(_T_981) + $signed(_T_977); // @[FixedPointTypeClass.scala 21:58]
  assign _T_984 = $signed(_T_983); // @[FixedPointTypeClass.scala 21:58]
  assign _T_986 = $signed(_T_984) + $signed(_T_978); // @[FixedPointTypeClass.scala 21:58]
  assign _T_987 = $signed(_T_986); // @[FixedPointTypeClass.scala 21:58]
  assign _T_988 = $signed(io_in_bits_0) * $signed(io_weightMatrix_76_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_989 = $signed(io_in_bits_1) * $signed(io_weightMatrix_76_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_990 = $signed(io_in_bits_2) * $signed(io_weightMatrix_76_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_991 = $signed(io_in_bits_3) * $signed(io_weightMatrix_76_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_993 = $signed(_T_988) + $signed(_T_989); // @[FixedPointTypeClass.scala 21:58]
  assign _T_994 = $signed(_T_993); // @[FixedPointTypeClass.scala 21:58]
  assign _T_996 = $signed(_T_994) + $signed(_T_990); // @[FixedPointTypeClass.scala 21:58]
  assign _T_997 = $signed(_T_996); // @[FixedPointTypeClass.scala 21:58]
  assign _T_999 = $signed(_T_997) + $signed(_T_991); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1000 = $signed(_T_999); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1001 = $signed(io_in_bits_0) * $signed(io_weightMatrix_77_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1002 = $signed(io_in_bits_1) * $signed(io_weightMatrix_77_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1003 = $signed(io_in_bits_2) * $signed(io_weightMatrix_77_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1004 = $signed(io_in_bits_3) * $signed(io_weightMatrix_77_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1006 = $signed(_T_1001) + $signed(_T_1002); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1007 = $signed(_T_1006); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1009 = $signed(_T_1007) + $signed(_T_1003); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1010 = $signed(_T_1009); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1012 = $signed(_T_1010) + $signed(_T_1004); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1013 = $signed(_T_1012); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1014 = $signed(io_in_bits_0) * $signed(io_weightMatrix_78_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1015 = $signed(io_in_bits_1) * $signed(io_weightMatrix_78_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1016 = $signed(io_in_bits_2) * $signed(io_weightMatrix_78_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1017 = $signed(io_in_bits_3) * $signed(io_weightMatrix_78_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1019 = $signed(_T_1014) + $signed(_T_1015); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1020 = $signed(_T_1019); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1022 = $signed(_T_1020) + $signed(_T_1016); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1023 = $signed(_T_1022); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1025 = $signed(_T_1023) + $signed(_T_1017); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1026 = $signed(_T_1025); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1027 = $signed(io_in_bits_0) * $signed(io_weightMatrix_79_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1028 = $signed(io_in_bits_1) * $signed(io_weightMatrix_79_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1029 = $signed(io_in_bits_2) * $signed(io_weightMatrix_79_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1030 = $signed(io_in_bits_3) * $signed(io_weightMatrix_79_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1032 = $signed(_T_1027) + $signed(_T_1028); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1033 = $signed(_T_1032); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1035 = $signed(_T_1033) + $signed(_T_1029); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1036 = $signed(_T_1035); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1038 = $signed(_T_1036) + $signed(_T_1030); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1039 = $signed(_T_1038); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1040 = $signed(io_in_bits_0) * $signed(io_weightMatrix_80_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1041 = $signed(io_in_bits_1) * $signed(io_weightMatrix_80_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1042 = $signed(io_in_bits_2) * $signed(io_weightMatrix_80_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1043 = $signed(io_in_bits_3) * $signed(io_weightMatrix_80_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1045 = $signed(_T_1040) + $signed(_T_1041); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1046 = $signed(_T_1045); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1048 = $signed(_T_1046) + $signed(_T_1042); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1049 = $signed(_T_1048); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1051 = $signed(_T_1049) + $signed(_T_1043); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1052 = $signed(_T_1051); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1053 = $signed(io_in_bits_0) * $signed(io_weightMatrix_81_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1054 = $signed(io_in_bits_1) * $signed(io_weightMatrix_81_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1055 = $signed(io_in_bits_2) * $signed(io_weightMatrix_81_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1056 = $signed(io_in_bits_3) * $signed(io_weightMatrix_81_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1058 = $signed(_T_1053) + $signed(_T_1054); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1059 = $signed(_T_1058); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1061 = $signed(_T_1059) + $signed(_T_1055); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1062 = $signed(_T_1061); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1064 = $signed(_T_1062) + $signed(_T_1056); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1065 = $signed(_T_1064); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1066 = $signed(io_in_bits_0) * $signed(io_weightMatrix_82_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1067 = $signed(io_in_bits_1) * $signed(io_weightMatrix_82_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1068 = $signed(io_in_bits_2) * $signed(io_weightMatrix_82_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1069 = $signed(io_in_bits_3) * $signed(io_weightMatrix_82_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1071 = $signed(_T_1066) + $signed(_T_1067); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1072 = $signed(_T_1071); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1074 = $signed(_T_1072) + $signed(_T_1068); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1075 = $signed(_T_1074); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1077 = $signed(_T_1075) + $signed(_T_1069); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1078 = $signed(_T_1077); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1079 = $signed(io_in_bits_0) * $signed(io_weightMatrix_83_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1080 = $signed(io_in_bits_1) * $signed(io_weightMatrix_83_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1081 = $signed(io_in_bits_2) * $signed(io_weightMatrix_83_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1082 = $signed(io_in_bits_3) * $signed(io_weightMatrix_83_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1084 = $signed(_T_1079) + $signed(_T_1080); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1085 = $signed(_T_1084); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1087 = $signed(_T_1085) + $signed(_T_1081); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1088 = $signed(_T_1087); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1090 = $signed(_T_1088) + $signed(_T_1082); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1091 = $signed(_T_1090); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1092 = $signed(io_in_bits_0) * $signed(io_weightMatrix_84_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1093 = $signed(io_in_bits_1) * $signed(io_weightMatrix_84_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1094 = $signed(io_in_bits_2) * $signed(io_weightMatrix_84_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1095 = $signed(io_in_bits_3) * $signed(io_weightMatrix_84_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1097 = $signed(_T_1092) + $signed(_T_1093); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1098 = $signed(_T_1097); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1100 = $signed(_T_1098) + $signed(_T_1094); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1101 = $signed(_T_1100); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1103 = $signed(_T_1101) + $signed(_T_1095); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1104 = $signed(_T_1103); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1105 = $signed(io_in_bits_0) * $signed(io_weightMatrix_85_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1106 = $signed(io_in_bits_1) * $signed(io_weightMatrix_85_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1107 = $signed(io_in_bits_2) * $signed(io_weightMatrix_85_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1108 = $signed(io_in_bits_3) * $signed(io_weightMatrix_85_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1110 = $signed(_T_1105) + $signed(_T_1106); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1111 = $signed(_T_1110); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1113 = $signed(_T_1111) + $signed(_T_1107); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1114 = $signed(_T_1113); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1116 = $signed(_T_1114) + $signed(_T_1108); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1117 = $signed(_T_1116); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1118 = $signed(io_in_bits_0) * $signed(io_weightMatrix_86_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1119 = $signed(io_in_bits_1) * $signed(io_weightMatrix_86_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1120 = $signed(io_in_bits_2) * $signed(io_weightMatrix_86_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1121 = $signed(io_in_bits_3) * $signed(io_weightMatrix_86_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1123 = $signed(_T_1118) + $signed(_T_1119); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1124 = $signed(_T_1123); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1126 = $signed(_T_1124) + $signed(_T_1120); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1127 = $signed(_T_1126); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1129 = $signed(_T_1127) + $signed(_T_1121); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1130 = $signed(_T_1129); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1131 = $signed(io_in_bits_0) * $signed(io_weightMatrix_87_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1132 = $signed(io_in_bits_1) * $signed(io_weightMatrix_87_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1133 = $signed(io_in_bits_2) * $signed(io_weightMatrix_87_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1134 = $signed(io_in_bits_3) * $signed(io_weightMatrix_87_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1136 = $signed(_T_1131) + $signed(_T_1132); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1137 = $signed(_T_1136); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1139 = $signed(_T_1137) + $signed(_T_1133); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1140 = $signed(_T_1139); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1142 = $signed(_T_1140) + $signed(_T_1134); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1143 = $signed(_T_1142); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1144 = $signed(io_in_bits_0) * $signed(io_weightMatrix_88_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1145 = $signed(io_in_bits_1) * $signed(io_weightMatrix_88_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1146 = $signed(io_in_bits_2) * $signed(io_weightMatrix_88_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1147 = $signed(io_in_bits_3) * $signed(io_weightMatrix_88_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1149 = $signed(_T_1144) + $signed(_T_1145); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1150 = $signed(_T_1149); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1152 = $signed(_T_1150) + $signed(_T_1146); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1153 = $signed(_T_1152); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1155 = $signed(_T_1153) + $signed(_T_1147); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1156 = $signed(_T_1155); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1157 = $signed(io_in_bits_0) * $signed(io_weightMatrix_89_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1158 = $signed(io_in_bits_1) * $signed(io_weightMatrix_89_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1159 = $signed(io_in_bits_2) * $signed(io_weightMatrix_89_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1160 = $signed(io_in_bits_3) * $signed(io_weightMatrix_89_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1162 = $signed(_T_1157) + $signed(_T_1158); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1163 = $signed(_T_1162); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1165 = $signed(_T_1163) + $signed(_T_1159); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1166 = $signed(_T_1165); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1168 = $signed(_T_1166) + $signed(_T_1160); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1169 = $signed(_T_1168); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1170 = $signed(io_in_bits_0) * $signed(io_weightMatrix_90_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1171 = $signed(io_in_bits_1) * $signed(io_weightMatrix_90_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1172 = $signed(io_in_bits_2) * $signed(io_weightMatrix_90_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1173 = $signed(io_in_bits_3) * $signed(io_weightMatrix_90_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1175 = $signed(_T_1170) + $signed(_T_1171); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1176 = $signed(_T_1175); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1178 = $signed(_T_1176) + $signed(_T_1172); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1179 = $signed(_T_1178); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1181 = $signed(_T_1179) + $signed(_T_1173); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1182 = $signed(_T_1181); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1183 = $signed(io_in_bits_0) * $signed(io_weightMatrix_91_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1184 = $signed(io_in_bits_1) * $signed(io_weightMatrix_91_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1185 = $signed(io_in_bits_2) * $signed(io_weightMatrix_91_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1186 = $signed(io_in_bits_3) * $signed(io_weightMatrix_91_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1188 = $signed(_T_1183) + $signed(_T_1184); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1189 = $signed(_T_1188); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1191 = $signed(_T_1189) + $signed(_T_1185); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1192 = $signed(_T_1191); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1194 = $signed(_T_1192) + $signed(_T_1186); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1195 = $signed(_T_1194); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1196 = $signed(io_in_bits_0) * $signed(io_weightMatrix_92_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1197 = $signed(io_in_bits_1) * $signed(io_weightMatrix_92_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1198 = $signed(io_in_bits_2) * $signed(io_weightMatrix_92_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1199 = $signed(io_in_bits_3) * $signed(io_weightMatrix_92_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1201 = $signed(_T_1196) + $signed(_T_1197); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1202 = $signed(_T_1201); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1204 = $signed(_T_1202) + $signed(_T_1198); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1205 = $signed(_T_1204); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1207 = $signed(_T_1205) + $signed(_T_1199); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1208 = $signed(_T_1207); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1209 = $signed(io_in_bits_0) * $signed(io_weightMatrix_93_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1210 = $signed(io_in_bits_1) * $signed(io_weightMatrix_93_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1211 = $signed(io_in_bits_2) * $signed(io_weightMatrix_93_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1212 = $signed(io_in_bits_3) * $signed(io_weightMatrix_93_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1214 = $signed(_T_1209) + $signed(_T_1210); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1215 = $signed(_T_1214); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1217 = $signed(_T_1215) + $signed(_T_1211); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1218 = $signed(_T_1217); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1220 = $signed(_T_1218) + $signed(_T_1212); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1221 = $signed(_T_1220); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1222 = $signed(io_in_bits_0) * $signed(io_weightMatrix_94_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1223 = $signed(io_in_bits_1) * $signed(io_weightMatrix_94_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1224 = $signed(io_in_bits_2) * $signed(io_weightMatrix_94_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1225 = $signed(io_in_bits_3) * $signed(io_weightMatrix_94_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1227 = $signed(_T_1222) + $signed(_T_1223); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1228 = $signed(_T_1227); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1230 = $signed(_T_1228) + $signed(_T_1224); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1231 = $signed(_T_1230); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1233 = $signed(_T_1231) + $signed(_T_1225); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1234 = $signed(_T_1233); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1235 = $signed(io_in_bits_0) * $signed(io_weightMatrix_95_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1236 = $signed(io_in_bits_1) * $signed(io_weightMatrix_95_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1237 = $signed(io_in_bits_2) * $signed(io_weightMatrix_95_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1238 = $signed(io_in_bits_3) * $signed(io_weightMatrix_95_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1240 = $signed(_T_1235) + $signed(_T_1236); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1241 = $signed(_T_1240); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1243 = $signed(_T_1241) + $signed(_T_1237); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1244 = $signed(_T_1243); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1246 = $signed(_T_1244) + $signed(_T_1238); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1247 = $signed(_T_1246); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1248 = $signed(io_in_bits_0) * $signed(io_weightMatrix_96_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1249 = $signed(io_in_bits_1) * $signed(io_weightMatrix_96_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1250 = $signed(io_in_bits_2) * $signed(io_weightMatrix_96_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1251 = $signed(io_in_bits_3) * $signed(io_weightMatrix_96_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1253 = $signed(_T_1248) + $signed(_T_1249); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1254 = $signed(_T_1253); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1256 = $signed(_T_1254) + $signed(_T_1250); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1257 = $signed(_T_1256); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1259 = $signed(_T_1257) + $signed(_T_1251); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1260 = $signed(_T_1259); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1261 = $signed(io_in_bits_0) * $signed(io_weightMatrix_97_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1262 = $signed(io_in_bits_1) * $signed(io_weightMatrix_97_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1263 = $signed(io_in_bits_2) * $signed(io_weightMatrix_97_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1264 = $signed(io_in_bits_3) * $signed(io_weightMatrix_97_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1266 = $signed(_T_1261) + $signed(_T_1262); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1267 = $signed(_T_1266); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1269 = $signed(_T_1267) + $signed(_T_1263); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1270 = $signed(_T_1269); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1272 = $signed(_T_1270) + $signed(_T_1264); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1273 = $signed(_T_1272); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1274 = $signed(io_in_bits_0) * $signed(io_weightMatrix_98_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1275 = $signed(io_in_bits_1) * $signed(io_weightMatrix_98_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1276 = $signed(io_in_bits_2) * $signed(io_weightMatrix_98_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1277 = $signed(io_in_bits_3) * $signed(io_weightMatrix_98_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1279 = $signed(_T_1274) + $signed(_T_1275); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1280 = $signed(_T_1279); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1282 = $signed(_T_1280) + $signed(_T_1276); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1283 = $signed(_T_1282); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1285 = $signed(_T_1283) + $signed(_T_1277); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1286 = $signed(_T_1285); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1287 = $signed(io_in_bits_0) * $signed(io_weightMatrix_99_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1288 = $signed(io_in_bits_1) * $signed(io_weightMatrix_99_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1289 = $signed(io_in_bits_2) * $signed(io_weightMatrix_99_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1290 = $signed(io_in_bits_3) * $signed(io_weightMatrix_99_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1292 = $signed(_T_1287) + $signed(_T_1288); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1293 = $signed(_T_1292); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1295 = $signed(_T_1293) + $signed(_T_1289); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1296 = $signed(_T_1295); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1298 = $signed(_T_1296) + $signed(_T_1290); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1299 = $signed(_T_1298); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_2 = _T_12[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_3 = _GEN_2[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_0 = $signed(_GEN_3); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1301 = $signed(inputWeighted_0) + $signed(io_biasVec_0); // @[FixedPointTypeClass.scala 21:58]
  assign biased_0 = $signed(_T_1301); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_4 = _T_25[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_5 = _GEN_4[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_1 = $signed(_GEN_5); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1304 = $signed(inputWeighted_1) + $signed(io_biasVec_1); // @[FixedPointTypeClass.scala 21:58]
  assign biased_1 = $signed(_T_1304); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_6 = _T_38[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_7 = _GEN_6[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_2 = $signed(_GEN_7); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1307 = $signed(inputWeighted_2) + $signed(io_biasVec_2); // @[FixedPointTypeClass.scala 21:58]
  assign biased_2 = $signed(_T_1307); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_8 = _T_51[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_9 = _GEN_8[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_3 = $signed(_GEN_9); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1310 = $signed(inputWeighted_3) + $signed(io_biasVec_3); // @[FixedPointTypeClass.scala 21:58]
  assign biased_3 = $signed(_T_1310); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_10 = _T_64[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_11 = _GEN_10[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_4 = $signed(_GEN_11); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1313 = $signed(inputWeighted_4) + $signed(io_biasVec_4); // @[FixedPointTypeClass.scala 21:58]
  assign biased_4 = $signed(_T_1313); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_12 = _T_77[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_13 = _GEN_12[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_5 = $signed(_GEN_13); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1316 = $signed(inputWeighted_5) + $signed(io_biasVec_5); // @[FixedPointTypeClass.scala 21:58]
  assign biased_5 = $signed(_T_1316); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_14 = _T_90[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_15 = _GEN_14[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_6 = $signed(_GEN_15); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1319 = $signed(inputWeighted_6) + $signed(io_biasVec_6); // @[FixedPointTypeClass.scala 21:58]
  assign biased_6 = $signed(_T_1319); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_16 = _T_103[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_17 = _GEN_16[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_7 = $signed(_GEN_17); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1322 = $signed(inputWeighted_7) + $signed(io_biasVec_7); // @[FixedPointTypeClass.scala 21:58]
  assign biased_7 = $signed(_T_1322); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_18 = _T_116[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_19 = _GEN_18[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_8 = $signed(_GEN_19); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1325 = $signed(inputWeighted_8) + $signed(io_biasVec_8); // @[FixedPointTypeClass.scala 21:58]
  assign biased_8 = $signed(_T_1325); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_20 = _T_129[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_21 = _GEN_20[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_9 = $signed(_GEN_21); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1328 = $signed(inputWeighted_9) + $signed(io_biasVec_9); // @[FixedPointTypeClass.scala 21:58]
  assign biased_9 = $signed(_T_1328); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_22 = _T_142[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_23 = _GEN_22[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_10 = $signed(_GEN_23); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1331 = $signed(inputWeighted_10) + $signed(io_biasVec_10); // @[FixedPointTypeClass.scala 21:58]
  assign biased_10 = $signed(_T_1331); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_24 = _T_155[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_25 = _GEN_24[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_11 = $signed(_GEN_25); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1334 = $signed(inputWeighted_11) + $signed(io_biasVec_11); // @[FixedPointTypeClass.scala 21:58]
  assign biased_11 = $signed(_T_1334); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_26 = _T_168[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_27 = _GEN_26[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_12 = $signed(_GEN_27); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1337 = $signed(inputWeighted_12) + $signed(io_biasVec_12); // @[FixedPointTypeClass.scala 21:58]
  assign biased_12 = $signed(_T_1337); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_28 = _T_181[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_29 = _GEN_28[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_13 = $signed(_GEN_29); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1340 = $signed(inputWeighted_13) + $signed(io_biasVec_13); // @[FixedPointTypeClass.scala 21:58]
  assign biased_13 = $signed(_T_1340); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_30 = _T_194[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_31 = _GEN_30[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_14 = $signed(_GEN_31); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1343 = $signed(inputWeighted_14) + $signed(io_biasVec_14); // @[FixedPointTypeClass.scala 21:58]
  assign biased_14 = $signed(_T_1343); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_32 = _T_207[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_33 = _GEN_32[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_15 = $signed(_GEN_33); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1346 = $signed(inputWeighted_15) + $signed(io_biasVec_15); // @[FixedPointTypeClass.scala 21:58]
  assign biased_15 = $signed(_T_1346); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_34 = _T_220[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_35 = _GEN_34[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_16 = $signed(_GEN_35); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1349 = $signed(inputWeighted_16) + $signed(io_biasVec_16); // @[FixedPointTypeClass.scala 21:58]
  assign biased_16 = $signed(_T_1349); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_36 = _T_233[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_37 = _GEN_36[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_17 = $signed(_GEN_37); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1352 = $signed(inputWeighted_17) + $signed(io_biasVec_17); // @[FixedPointTypeClass.scala 21:58]
  assign biased_17 = $signed(_T_1352); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_38 = _T_246[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_39 = _GEN_38[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_18 = $signed(_GEN_39); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1355 = $signed(inputWeighted_18) + $signed(io_biasVec_18); // @[FixedPointTypeClass.scala 21:58]
  assign biased_18 = $signed(_T_1355); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_40 = _T_259[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_41 = _GEN_40[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_19 = $signed(_GEN_41); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1358 = $signed(inputWeighted_19) + $signed(io_biasVec_19); // @[FixedPointTypeClass.scala 21:58]
  assign biased_19 = $signed(_T_1358); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_42 = _T_272[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_43 = _GEN_42[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_20 = $signed(_GEN_43); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1361 = $signed(inputWeighted_20) + $signed(io_biasVec_20); // @[FixedPointTypeClass.scala 21:58]
  assign biased_20 = $signed(_T_1361); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_44 = _T_285[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_45 = _GEN_44[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_21 = $signed(_GEN_45); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1364 = $signed(inputWeighted_21) + $signed(io_biasVec_21); // @[FixedPointTypeClass.scala 21:58]
  assign biased_21 = $signed(_T_1364); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_46 = _T_298[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_47 = _GEN_46[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_22 = $signed(_GEN_47); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1367 = $signed(inputWeighted_22) + $signed(io_biasVec_22); // @[FixedPointTypeClass.scala 21:58]
  assign biased_22 = $signed(_T_1367); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_48 = _T_311[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_49 = _GEN_48[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_23 = $signed(_GEN_49); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1370 = $signed(inputWeighted_23) + $signed(io_biasVec_23); // @[FixedPointTypeClass.scala 21:58]
  assign biased_23 = $signed(_T_1370); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_50 = _T_324[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_51 = _GEN_50[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_24 = $signed(_GEN_51); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1373 = $signed(inputWeighted_24) + $signed(io_biasVec_24); // @[FixedPointTypeClass.scala 21:58]
  assign biased_24 = $signed(_T_1373); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_52 = _T_337[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_53 = _GEN_52[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_25 = $signed(_GEN_53); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1376 = $signed(inputWeighted_25) + $signed(io_biasVec_25); // @[FixedPointTypeClass.scala 21:58]
  assign biased_25 = $signed(_T_1376); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_54 = _T_350[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_55 = _GEN_54[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_26 = $signed(_GEN_55); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1379 = $signed(inputWeighted_26) + $signed(io_biasVec_26); // @[FixedPointTypeClass.scala 21:58]
  assign biased_26 = $signed(_T_1379); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_56 = _T_363[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_57 = _GEN_56[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_27 = $signed(_GEN_57); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1382 = $signed(inputWeighted_27) + $signed(io_biasVec_27); // @[FixedPointTypeClass.scala 21:58]
  assign biased_27 = $signed(_T_1382); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_58 = _T_376[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_59 = _GEN_58[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_28 = $signed(_GEN_59); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1385 = $signed(inputWeighted_28) + $signed(io_biasVec_28); // @[FixedPointTypeClass.scala 21:58]
  assign biased_28 = $signed(_T_1385); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_60 = _T_389[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_61 = _GEN_60[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_29 = $signed(_GEN_61); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1388 = $signed(inputWeighted_29) + $signed(io_biasVec_29); // @[FixedPointTypeClass.scala 21:58]
  assign biased_29 = $signed(_T_1388); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_62 = _T_402[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_63 = _GEN_62[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_30 = $signed(_GEN_63); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1391 = $signed(inputWeighted_30) + $signed(io_biasVec_30); // @[FixedPointTypeClass.scala 21:58]
  assign biased_30 = $signed(_T_1391); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_64 = _T_415[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_65 = _GEN_64[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_31 = $signed(_GEN_65); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1394 = $signed(inputWeighted_31) + $signed(io_biasVec_31); // @[FixedPointTypeClass.scala 21:58]
  assign biased_31 = $signed(_T_1394); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_66 = _T_428[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_67 = _GEN_66[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_32 = $signed(_GEN_67); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1397 = $signed(inputWeighted_32) + $signed(io_biasVec_32); // @[FixedPointTypeClass.scala 21:58]
  assign biased_32 = $signed(_T_1397); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_68 = _T_441[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_69 = _GEN_68[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_33 = $signed(_GEN_69); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1400 = $signed(inputWeighted_33) + $signed(io_biasVec_33); // @[FixedPointTypeClass.scala 21:58]
  assign biased_33 = $signed(_T_1400); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_70 = _T_454[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_71 = _GEN_70[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_34 = $signed(_GEN_71); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1403 = $signed(inputWeighted_34) + $signed(io_biasVec_34); // @[FixedPointTypeClass.scala 21:58]
  assign biased_34 = $signed(_T_1403); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_72 = _T_467[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_73 = _GEN_72[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_35 = $signed(_GEN_73); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1406 = $signed(inputWeighted_35) + $signed(io_biasVec_35); // @[FixedPointTypeClass.scala 21:58]
  assign biased_35 = $signed(_T_1406); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_74 = _T_480[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_75 = _GEN_74[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_36 = $signed(_GEN_75); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1409 = $signed(inputWeighted_36) + $signed(io_biasVec_36); // @[FixedPointTypeClass.scala 21:58]
  assign biased_36 = $signed(_T_1409); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_76 = _T_493[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_77 = _GEN_76[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_37 = $signed(_GEN_77); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1412 = $signed(inputWeighted_37) + $signed(io_biasVec_37); // @[FixedPointTypeClass.scala 21:58]
  assign biased_37 = $signed(_T_1412); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_78 = _T_506[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_79 = _GEN_78[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_38 = $signed(_GEN_79); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1415 = $signed(inputWeighted_38) + $signed(io_biasVec_38); // @[FixedPointTypeClass.scala 21:58]
  assign biased_38 = $signed(_T_1415); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_80 = _T_519[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_81 = _GEN_80[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_39 = $signed(_GEN_81); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1418 = $signed(inputWeighted_39) + $signed(io_biasVec_39); // @[FixedPointTypeClass.scala 21:58]
  assign biased_39 = $signed(_T_1418); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_82 = _T_532[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_83 = _GEN_82[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_40 = $signed(_GEN_83); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1421 = $signed(inputWeighted_40) + $signed(io_biasVec_40); // @[FixedPointTypeClass.scala 21:58]
  assign biased_40 = $signed(_T_1421); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_84 = _T_545[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_85 = _GEN_84[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_41 = $signed(_GEN_85); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1424 = $signed(inputWeighted_41) + $signed(io_biasVec_41); // @[FixedPointTypeClass.scala 21:58]
  assign biased_41 = $signed(_T_1424); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_86 = _T_558[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_87 = _GEN_86[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_42 = $signed(_GEN_87); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1427 = $signed(inputWeighted_42) + $signed(io_biasVec_42); // @[FixedPointTypeClass.scala 21:58]
  assign biased_42 = $signed(_T_1427); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_88 = _T_571[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_89 = _GEN_88[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_43 = $signed(_GEN_89); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1430 = $signed(inputWeighted_43) + $signed(io_biasVec_43); // @[FixedPointTypeClass.scala 21:58]
  assign biased_43 = $signed(_T_1430); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_90 = _T_584[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_91 = _GEN_90[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_44 = $signed(_GEN_91); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1433 = $signed(inputWeighted_44) + $signed(io_biasVec_44); // @[FixedPointTypeClass.scala 21:58]
  assign biased_44 = $signed(_T_1433); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_92 = _T_597[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_93 = _GEN_92[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_45 = $signed(_GEN_93); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1436 = $signed(inputWeighted_45) + $signed(io_biasVec_45); // @[FixedPointTypeClass.scala 21:58]
  assign biased_45 = $signed(_T_1436); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_94 = _T_610[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_95 = _GEN_94[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_46 = $signed(_GEN_95); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1439 = $signed(inputWeighted_46) + $signed(io_biasVec_46); // @[FixedPointTypeClass.scala 21:58]
  assign biased_46 = $signed(_T_1439); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_96 = _T_623[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_97 = _GEN_96[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_47 = $signed(_GEN_97); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1442 = $signed(inputWeighted_47) + $signed(io_biasVec_47); // @[FixedPointTypeClass.scala 21:58]
  assign biased_47 = $signed(_T_1442); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_98 = _T_636[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_99 = _GEN_98[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_48 = $signed(_GEN_99); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1445 = $signed(inputWeighted_48) + $signed(io_biasVec_48); // @[FixedPointTypeClass.scala 21:58]
  assign biased_48 = $signed(_T_1445); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_100 = _T_649[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_101 = _GEN_100[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_49 = $signed(_GEN_101); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1448 = $signed(inputWeighted_49) + $signed(io_biasVec_49); // @[FixedPointTypeClass.scala 21:58]
  assign biased_49 = $signed(_T_1448); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_102 = _T_662[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_103 = _GEN_102[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_50 = $signed(_GEN_103); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1451 = $signed(inputWeighted_50) + $signed(io_biasVec_50); // @[FixedPointTypeClass.scala 21:58]
  assign biased_50 = $signed(_T_1451); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_104 = _T_675[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_105 = _GEN_104[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_51 = $signed(_GEN_105); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1454 = $signed(inputWeighted_51) + $signed(io_biasVec_51); // @[FixedPointTypeClass.scala 21:58]
  assign biased_51 = $signed(_T_1454); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_106 = _T_688[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_107 = _GEN_106[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_52 = $signed(_GEN_107); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1457 = $signed(inputWeighted_52) + $signed(io_biasVec_52); // @[FixedPointTypeClass.scala 21:58]
  assign biased_52 = $signed(_T_1457); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_108 = _T_701[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_109 = _GEN_108[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_53 = $signed(_GEN_109); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1460 = $signed(inputWeighted_53) + $signed(io_biasVec_53); // @[FixedPointTypeClass.scala 21:58]
  assign biased_53 = $signed(_T_1460); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_110 = _T_714[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_111 = _GEN_110[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_54 = $signed(_GEN_111); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1463 = $signed(inputWeighted_54) + $signed(io_biasVec_54); // @[FixedPointTypeClass.scala 21:58]
  assign biased_54 = $signed(_T_1463); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_112 = _T_727[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_113 = _GEN_112[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_55 = $signed(_GEN_113); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1466 = $signed(inputWeighted_55) + $signed(io_biasVec_55); // @[FixedPointTypeClass.scala 21:58]
  assign biased_55 = $signed(_T_1466); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_114 = _T_740[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_115 = _GEN_114[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_56 = $signed(_GEN_115); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1469 = $signed(inputWeighted_56) + $signed(io_biasVec_56); // @[FixedPointTypeClass.scala 21:58]
  assign biased_56 = $signed(_T_1469); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_116 = _T_753[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_117 = _GEN_116[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_57 = $signed(_GEN_117); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1472 = $signed(inputWeighted_57) + $signed(io_biasVec_57); // @[FixedPointTypeClass.scala 21:58]
  assign biased_57 = $signed(_T_1472); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_118 = _T_766[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_119 = _GEN_118[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_58 = $signed(_GEN_119); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1475 = $signed(inputWeighted_58) + $signed(io_biasVec_58); // @[FixedPointTypeClass.scala 21:58]
  assign biased_58 = $signed(_T_1475); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_120 = _T_779[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_121 = _GEN_120[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_59 = $signed(_GEN_121); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1478 = $signed(inputWeighted_59) + $signed(io_biasVec_59); // @[FixedPointTypeClass.scala 21:58]
  assign biased_59 = $signed(_T_1478); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_122 = _T_792[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_123 = _GEN_122[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_60 = $signed(_GEN_123); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1481 = $signed(inputWeighted_60) + $signed(io_biasVec_60); // @[FixedPointTypeClass.scala 21:58]
  assign biased_60 = $signed(_T_1481); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_124 = _T_805[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_125 = _GEN_124[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_61 = $signed(_GEN_125); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1484 = $signed(inputWeighted_61) + $signed(io_biasVec_61); // @[FixedPointTypeClass.scala 21:58]
  assign biased_61 = $signed(_T_1484); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_126 = _T_818[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_127 = _GEN_126[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_62 = $signed(_GEN_127); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1487 = $signed(inputWeighted_62) + $signed(io_biasVec_62); // @[FixedPointTypeClass.scala 21:58]
  assign biased_62 = $signed(_T_1487); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_128 = _T_831[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_129 = _GEN_128[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_63 = $signed(_GEN_129); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1490 = $signed(inputWeighted_63) + $signed(io_biasVec_63); // @[FixedPointTypeClass.scala 21:58]
  assign biased_63 = $signed(_T_1490); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_130 = _T_844[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_131 = _GEN_130[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_64 = $signed(_GEN_131); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1493 = $signed(inputWeighted_64) + $signed(io_biasVec_64); // @[FixedPointTypeClass.scala 21:58]
  assign biased_64 = $signed(_T_1493); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_132 = _T_857[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_133 = _GEN_132[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_65 = $signed(_GEN_133); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1496 = $signed(inputWeighted_65) + $signed(io_biasVec_65); // @[FixedPointTypeClass.scala 21:58]
  assign biased_65 = $signed(_T_1496); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_134 = _T_870[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_135 = _GEN_134[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_66 = $signed(_GEN_135); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1499 = $signed(inputWeighted_66) + $signed(io_biasVec_66); // @[FixedPointTypeClass.scala 21:58]
  assign biased_66 = $signed(_T_1499); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_136 = _T_883[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_137 = _GEN_136[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_67 = $signed(_GEN_137); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1502 = $signed(inputWeighted_67) + $signed(io_biasVec_67); // @[FixedPointTypeClass.scala 21:58]
  assign biased_67 = $signed(_T_1502); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_138 = _T_896[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_139 = _GEN_138[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_68 = $signed(_GEN_139); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1505 = $signed(inputWeighted_68) + $signed(io_biasVec_68); // @[FixedPointTypeClass.scala 21:58]
  assign biased_68 = $signed(_T_1505); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_140 = _T_909[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_141 = _GEN_140[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_69 = $signed(_GEN_141); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1508 = $signed(inputWeighted_69) + $signed(io_biasVec_69); // @[FixedPointTypeClass.scala 21:58]
  assign biased_69 = $signed(_T_1508); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_142 = _T_922[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_143 = _GEN_142[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_70 = $signed(_GEN_143); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1511 = $signed(inputWeighted_70) + $signed(io_biasVec_70); // @[FixedPointTypeClass.scala 21:58]
  assign biased_70 = $signed(_T_1511); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_144 = _T_935[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_145 = _GEN_144[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_71 = $signed(_GEN_145); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1514 = $signed(inputWeighted_71) + $signed(io_biasVec_71); // @[FixedPointTypeClass.scala 21:58]
  assign biased_71 = $signed(_T_1514); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_146 = _T_948[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_147 = _GEN_146[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_72 = $signed(_GEN_147); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1517 = $signed(inputWeighted_72) + $signed(io_biasVec_72); // @[FixedPointTypeClass.scala 21:58]
  assign biased_72 = $signed(_T_1517); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_148 = _T_961[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_149 = _GEN_148[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_73 = $signed(_GEN_149); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1520 = $signed(inputWeighted_73) + $signed(io_biasVec_73); // @[FixedPointTypeClass.scala 21:58]
  assign biased_73 = $signed(_T_1520); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_150 = _T_974[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_151 = _GEN_150[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_74 = $signed(_GEN_151); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1523 = $signed(inputWeighted_74) + $signed(io_biasVec_74); // @[FixedPointTypeClass.scala 21:58]
  assign biased_74 = $signed(_T_1523); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_152 = _T_987[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_153 = _GEN_152[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_75 = $signed(_GEN_153); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1526 = $signed(inputWeighted_75) + $signed(io_biasVec_75); // @[FixedPointTypeClass.scala 21:58]
  assign biased_75 = $signed(_T_1526); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_154 = _T_1000[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_155 = _GEN_154[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_76 = $signed(_GEN_155); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1529 = $signed(inputWeighted_76) + $signed(io_biasVec_76); // @[FixedPointTypeClass.scala 21:58]
  assign biased_76 = $signed(_T_1529); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_156 = _T_1013[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_157 = _GEN_156[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_77 = $signed(_GEN_157); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1532 = $signed(inputWeighted_77) + $signed(io_biasVec_77); // @[FixedPointTypeClass.scala 21:58]
  assign biased_77 = $signed(_T_1532); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_158 = _T_1026[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_159 = _GEN_158[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_78 = $signed(_GEN_159); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1535 = $signed(inputWeighted_78) + $signed(io_biasVec_78); // @[FixedPointTypeClass.scala 21:58]
  assign biased_78 = $signed(_T_1535); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_160 = _T_1039[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_161 = _GEN_160[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_79 = $signed(_GEN_161); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1538 = $signed(inputWeighted_79) + $signed(io_biasVec_79); // @[FixedPointTypeClass.scala 21:58]
  assign biased_79 = $signed(_T_1538); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_162 = _T_1052[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_163 = _GEN_162[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_80 = $signed(_GEN_163); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1541 = $signed(inputWeighted_80) + $signed(io_biasVec_80); // @[FixedPointTypeClass.scala 21:58]
  assign biased_80 = $signed(_T_1541); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_164 = _T_1065[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_165 = _GEN_164[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_81 = $signed(_GEN_165); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1544 = $signed(inputWeighted_81) + $signed(io_biasVec_81); // @[FixedPointTypeClass.scala 21:58]
  assign biased_81 = $signed(_T_1544); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_166 = _T_1078[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_167 = _GEN_166[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_82 = $signed(_GEN_167); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1547 = $signed(inputWeighted_82) + $signed(io_biasVec_82); // @[FixedPointTypeClass.scala 21:58]
  assign biased_82 = $signed(_T_1547); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_168 = _T_1091[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_169 = _GEN_168[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_83 = $signed(_GEN_169); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1550 = $signed(inputWeighted_83) + $signed(io_biasVec_83); // @[FixedPointTypeClass.scala 21:58]
  assign biased_83 = $signed(_T_1550); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_170 = _T_1104[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_171 = _GEN_170[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_84 = $signed(_GEN_171); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1553 = $signed(inputWeighted_84) + $signed(io_biasVec_84); // @[FixedPointTypeClass.scala 21:58]
  assign biased_84 = $signed(_T_1553); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_172 = _T_1117[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_173 = _GEN_172[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_85 = $signed(_GEN_173); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1556 = $signed(inputWeighted_85) + $signed(io_biasVec_85); // @[FixedPointTypeClass.scala 21:58]
  assign biased_85 = $signed(_T_1556); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_174 = _T_1130[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_175 = _GEN_174[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_86 = $signed(_GEN_175); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1559 = $signed(inputWeighted_86) + $signed(io_biasVec_86); // @[FixedPointTypeClass.scala 21:58]
  assign biased_86 = $signed(_T_1559); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_176 = _T_1143[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_177 = _GEN_176[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_87 = $signed(_GEN_177); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1562 = $signed(inputWeighted_87) + $signed(io_biasVec_87); // @[FixedPointTypeClass.scala 21:58]
  assign biased_87 = $signed(_T_1562); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_178 = _T_1156[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_179 = _GEN_178[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_88 = $signed(_GEN_179); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1565 = $signed(inputWeighted_88) + $signed(io_biasVec_88); // @[FixedPointTypeClass.scala 21:58]
  assign biased_88 = $signed(_T_1565); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_180 = _T_1169[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_181 = _GEN_180[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_89 = $signed(_GEN_181); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1568 = $signed(inputWeighted_89) + $signed(io_biasVec_89); // @[FixedPointTypeClass.scala 21:58]
  assign biased_89 = $signed(_T_1568); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_182 = _T_1182[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_183 = _GEN_182[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_90 = $signed(_GEN_183); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1571 = $signed(inputWeighted_90) + $signed(io_biasVec_90); // @[FixedPointTypeClass.scala 21:58]
  assign biased_90 = $signed(_T_1571); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_184 = _T_1195[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_185 = _GEN_184[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_91 = $signed(_GEN_185); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1574 = $signed(inputWeighted_91) + $signed(io_biasVec_91); // @[FixedPointTypeClass.scala 21:58]
  assign biased_91 = $signed(_T_1574); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_186 = _T_1208[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_187 = _GEN_186[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_92 = $signed(_GEN_187); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1577 = $signed(inputWeighted_92) + $signed(io_biasVec_92); // @[FixedPointTypeClass.scala 21:58]
  assign biased_92 = $signed(_T_1577); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_188 = _T_1221[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_189 = _GEN_188[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_93 = $signed(_GEN_189); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1580 = $signed(inputWeighted_93) + $signed(io_biasVec_93); // @[FixedPointTypeClass.scala 21:58]
  assign biased_93 = $signed(_T_1580); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_190 = _T_1234[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_191 = _GEN_190[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_94 = $signed(_GEN_191); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1583 = $signed(inputWeighted_94) + $signed(io_biasVec_94); // @[FixedPointTypeClass.scala 21:58]
  assign biased_94 = $signed(_T_1583); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_192 = _T_1247[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_193 = _GEN_192[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_95 = $signed(_GEN_193); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1586 = $signed(inputWeighted_95) + $signed(io_biasVec_95); // @[FixedPointTypeClass.scala 21:58]
  assign biased_95 = $signed(_T_1586); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_194 = _T_1260[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_195 = _GEN_194[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_96 = $signed(_GEN_195); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1589 = $signed(inputWeighted_96) + $signed(io_biasVec_96); // @[FixedPointTypeClass.scala 21:58]
  assign biased_96 = $signed(_T_1589); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_196 = _T_1273[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_197 = _GEN_196[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_97 = $signed(_GEN_197); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1592 = $signed(inputWeighted_97) + $signed(io_biasVec_97); // @[FixedPointTypeClass.scala 21:58]
  assign biased_97 = $signed(_T_1592); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_198 = _T_1286[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_199 = _GEN_198[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_98 = $signed(_GEN_199); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1595 = $signed(inputWeighted_98) + $signed(io_biasVec_98); // @[FixedPointTypeClass.scala 21:58]
  assign biased_98 = $signed(_T_1595); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_200 = _T_1299[63:8]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _GEN_201 = _GEN_200[31:0]; // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign inputWeighted_99 = $signed(_GEN_201); // @[neuralNet.scala 50:27 neuralNet.scala 52:22]
  assign _T_1598 = $signed(inputWeighted_99) + $signed(io_biasVec_99); // @[FixedPointTypeClass.scala 21:58]
  assign biased_99 = $signed(_T_1598); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1600 = $signed(biased_0) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_0 = _T_1600 ? $signed(biased_0) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1602 = $signed(biased_1) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_1 = _T_1602 ? $signed(biased_1) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1604 = $signed(biased_2) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_2 = _T_1604 ? $signed(biased_2) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1606 = $signed(biased_3) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_3 = _T_1606 ? $signed(biased_3) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1608 = $signed(biased_4) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_4 = _T_1608 ? $signed(biased_4) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1610 = $signed(biased_5) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_5 = _T_1610 ? $signed(biased_5) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1612 = $signed(biased_6) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_6 = _T_1612 ? $signed(biased_6) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1614 = $signed(biased_7) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_7 = _T_1614 ? $signed(biased_7) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1616 = $signed(biased_8) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_8 = _T_1616 ? $signed(biased_8) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1618 = $signed(biased_9) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_9 = _T_1618 ? $signed(biased_9) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1620 = $signed(biased_10) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_10 = _T_1620 ? $signed(biased_10) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1622 = $signed(biased_11) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_11 = _T_1622 ? $signed(biased_11) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1624 = $signed(biased_12) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_12 = _T_1624 ? $signed(biased_12) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1626 = $signed(biased_13) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_13 = _T_1626 ? $signed(biased_13) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1628 = $signed(biased_14) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_14 = _T_1628 ? $signed(biased_14) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1630 = $signed(biased_15) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_15 = _T_1630 ? $signed(biased_15) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1632 = $signed(biased_16) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_16 = _T_1632 ? $signed(biased_16) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1634 = $signed(biased_17) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_17 = _T_1634 ? $signed(biased_17) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1636 = $signed(biased_18) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_18 = _T_1636 ? $signed(biased_18) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1638 = $signed(biased_19) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_19 = _T_1638 ? $signed(biased_19) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1640 = $signed(biased_20) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_20 = _T_1640 ? $signed(biased_20) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1642 = $signed(biased_21) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_21 = _T_1642 ? $signed(biased_21) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1644 = $signed(biased_22) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_22 = _T_1644 ? $signed(biased_22) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1646 = $signed(biased_23) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_23 = _T_1646 ? $signed(biased_23) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1648 = $signed(biased_24) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_24 = _T_1648 ? $signed(biased_24) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1650 = $signed(biased_25) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_25 = _T_1650 ? $signed(biased_25) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1652 = $signed(biased_26) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_26 = _T_1652 ? $signed(biased_26) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1654 = $signed(biased_27) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_27 = _T_1654 ? $signed(biased_27) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1656 = $signed(biased_28) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_28 = _T_1656 ? $signed(biased_28) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1658 = $signed(biased_29) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_29 = _T_1658 ? $signed(biased_29) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1660 = $signed(biased_30) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_30 = _T_1660 ? $signed(biased_30) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1662 = $signed(biased_31) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_31 = _T_1662 ? $signed(biased_31) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1664 = $signed(biased_32) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_32 = _T_1664 ? $signed(biased_32) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1666 = $signed(biased_33) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_33 = _T_1666 ? $signed(biased_33) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1668 = $signed(biased_34) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_34 = _T_1668 ? $signed(biased_34) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1670 = $signed(biased_35) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_35 = _T_1670 ? $signed(biased_35) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1672 = $signed(biased_36) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_36 = _T_1672 ? $signed(biased_36) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1674 = $signed(biased_37) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_37 = _T_1674 ? $signed(biased_37) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1676 = $signed(biased_38) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_38 = _T_1676 ? $signed(biased_38) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1678 = $signed(biased_39) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_39 = _T_1678 ? $signed(biased_39) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1680 = $signed(biased_40) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_40 = _T_1680 ? $signed(biased_40) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1682 = $signed(biased_41) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_41 = _T_1682 ? $signed(biased_41) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1684 = $signed(biased_42) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_42 = _T_1684 ? $signed(biased_42) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1686 = $signed(biased_43) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_43 = _T_1686 ? $signed(biased_43) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1688 = $signed(biased_44) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_44 = _T_1688 ? $signed(biased_44) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1690 = $signed(biased_45) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_45 = _T_1690 ? $signed(biased_45) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1692 = $signed(biased_46) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_46 = _T_1692 ? $signed(biased_46) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1694 = $signed(biased_47) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_47 = _T_1694 ? $signed(biased_47) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1696 = $signed(biased_48) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_48 = _T_1696 ? $signed(biased_48) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1698 = $signed(biased_49) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_49 = _T_1698 ? $signed(biased_49) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1700 = $signed(biased_50) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_50 = _T_1700 ? $signed(biased_50) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1702 = $signed(biased_51) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_51 = _T_1702 ? $signed(biased_51) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1704 = $signed(biased_52) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_52 = _T_1704 ? $signed(biased_52) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1706 = $signed(biased_53) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_53 = _T_1706 ? $signed(biased_53) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1708 = $signed(biased_54) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_54 = _T_1708 ? $signed(biased_54) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1710 = $signed(biased_55) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_55 = _T_1710 ? $signed(biased_55) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1712 = $signed(biased_56) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_56 = _T_1712 ? $signed(biased_56) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1714 = $signed(biased_57) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_57 = _T_1714 ? $signed(biased_57) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1716 = $signed(biased_58) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_58 = _T_1716 ? $signed(biased_58) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1718 = $signed(biased_59) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_59 = _T_1718 ? $signed(biased_59) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1720 = $signed(biased_60) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_60 = _T_1720 ? $signed(biased_60) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1722 = $signed(biased_61) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_61 = _T_1722 ? $signed(biased_61) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1724 = $signed(biased_62) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_62 = _T_1724 ? $signed(biased_62) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1726 = $signed(biased_63) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_63 = _T_1726 ? $signed(biased_63) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1728 = $signed(biased_64) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_64 = _T_1728 ? $signed(biased_64) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1730 = $signed(biased_65) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_65 = _T_1730 ? $signed(biased_65) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1732 = $signed(biased_66) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_66 = _T_1732 ? $signed(biased_66) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1734 = $signed(biased_67) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_67 = _T_1734 ? $signed(biased_67) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1736 = $signed(biased_68) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_68 = _T_1736 ? $signed(biased_68) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1738 = $signed(biased_69) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_69 = _T_1738 ? $signed(biased_69) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1740 = $signed(biased_70) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_70 = _T_1740 ? $signed(biased_70) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1742 = $signed(biased_71) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_71 = _T_1742 ? $signed(biased_71) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1744 = $signed(biased_72) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_72 = _T_1744 ? $signed(biased_72) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1746 = $signed(biased_73) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_73 = _T_1746 ? $signed(biased_73) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1748 = $signed(biased_74) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_74 = _T_1748 ? $signed(biased_74) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1750 = $signed(biased_75) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_75 = _T_1750 ? $signed(biased_75) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1752 = $signed(biased_76) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_76 = _T_1752 ? $signed(biased_76) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1754 = $signed(biased_77) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_77 = _T_1754 ? $signed(biased_77) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1756 = $signed(biased_78) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_78 = _T_1756 ? $signed(biased_78) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1758 = $signed(biased_79) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_79 = _T_1758 ? $signed(biased_79) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1760 = $signed(biased_80) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_80 = _T_1760 ? $signed(biased_80) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1762 = $signed(biased_81) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_81 = _T_1762 ? $signed(biased_81) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1764 = $signed(biased_82) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_82 = _T_1764 ? $signed(biased_82) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1766 = $signed(biased_83) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_83 = _T_1766 ? $signed(biased_83) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1768 = $signed(biased_84) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_84 = _T_1768 ? $signed(biased_84) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1770 = $signed(biased_85) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_85 = _T_1770 ? $signed(biased_85) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1772 = $signed(biased_86) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_86 = _T_1772 ? $signed(biased_86) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1774 = $signed(biased_87) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_87 = _T_1774 ? $signed(biased_87) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1776 = $signed(biased_88) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_88 = _T_1776 ? $signed(biased_88) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1778 = $signed(biased_89) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_89 = _T_1778 ? $signed(biased_89) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1780 = $signed(biased_90) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_90 = _T_1780 ? $signed(biased_90) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1782 = $signed(biased_91) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_91 = _T_1782 ? $signed(biased_91) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1784 = $signed(biased_92) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_92 = _T_1784 ? $signed(biased_92) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1786 = $signed(biased_93) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_93 = _T_1786 ? $signed(biased_93) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1788 = $signed(biased_94) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_94 = _T_1788 ? $signed(biased_94) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1790 = $signed(biased_95) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_95 = _T_1790 ? $signed(biased_95) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1792 = $signed(biased_96) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_96 = _T_1792 ? $signed(biased_96) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1794 = $signed(biased_97) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_97 = _T_1794 ? $signed(biased_97) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1796 = $signed(biased_98) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_98 = _T_1796 ? $signed(biased_98) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1798 = $signed(biased_99) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign hiddenLayer_99 = _T_1798 ? $signed(biased_99) : $signed(32'sh0); // @[neuralNet.scala 62:26]
  assign _T_1800 = $signed(hiddenLayer_0) * $signed(io_weightVec_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1801 = $signed(hiddenLayer_1) * $signed(io_weightVec_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1802 = $signed(hiddenLayer_2) * $signed(io_weightVec_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1803 = $signed(hiddenLayer_3) * $signed(io_weightVec_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1804 = $signed(hiddenLayer_4) * $signed(io_weightVec_4); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1805 = $signed(hiddenLayer_5) * $signed(io_weightVec_5); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1806 = $signed(hiddenLayer_6) * $signed(io_weightVec_6); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1807 = $signed(hiddenLayer_7) * $signed(io_weightVec_7); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1808 = $signed(hiddenLayer_8) * $signed(io_weightVec_8); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1809 = $signed(hiddenLayer_9) * $signed(io_weightVec_9); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1810 = $signed(hiddenLayer_10) * $signed(io_weightVec_10); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1811 = $signed(hiddenLayer_11) * $signed(io_weightVec_11); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1812 = $signed(hiddenLayer_12) * $signed(io_weightVec_12); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1813 = $signed(hiddenLayer_13) * $signed(io_weightVec_13); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1814 = $signed(hiddenLayer_14) * $signed(io_weightVec_14); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1815 = $signed(hiddenLayer_15) * $signed(io_weightVec_15); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1816 = $signed(hiddenLayer_16) * $signed(io_weightVec_16); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1817 = $signed(hiddenLayer_17) * $signed(io_weightVec_17); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1818 = $signed(hiddenLayer_18) * $signed(io_weightVec_18); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1819 = $signed(hiddenLayer_19) * $signed(io_weightVec_19); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1820 = $signed(hiddenLayer_20) * $signed(io_weightVec_20); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1821 = $signed(hiddenLayer_21) * $signed(io_weightVec_21); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1822 = $signed(hiddenLayer_22) * $signed(io_weightVec_22); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1823 = $signed(hiddenLayer_23) * $signed(io_weightVec_23); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1824 = $signed(hiddenLayer_24) * $signed(io_weightVec_24); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1825 = $signed(hiddenLayer_25) * $signed(io_weightVec_25); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1826 = $signed(hiddenLayer_26) * $signed(io_weightVec_26); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1827 = $signed(hiddenLayer_27) * $signed(io_weightVec_27); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1828 = $signed(hiddenLayer_28) * $signed(io_weightVec_28); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1829 = $signed(hiddenLayer_29) * $signed(io_weightVec_29); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1830 = $signed(hiddenLayer_30) * $signed(io_weightVec_30); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1831 = $signed(hiddenLayer_31) * $signed(io_weightVec_31); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1832 = $signed(hiddenLayer_32) * $signed(io_weightVec_32); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1833 = $signed(hiddenLayer_33) * $signed(io_weightVec_33); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1834 = $signed(hiddenLayer_34) * $signed(io_weightVec_34); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1835 = $signed(hiddenLayer_35) * $signed(io_weightVec_35); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1836 = $signed(hiddenLayer_36) * $signed(io_weightVec_36); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1837 = $signed(hiddenLayer_37) * $signed(io_weightVec_37); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1838 = $signed(hiddenLayer_38) * $signed(io_weightVec_38); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1839 = $signed(hiddenLayer_39) * $signed(io_weightVec_39); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1840 = $signed(hiddenLayer_40) * $signed(io_weightVec_40); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1841 = $signed(hiddenLayer_41) * $signed(io_weightVec_41); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1842 = $signed(hiddenLayer_42) * $signed(io_weightVec_42); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1843 = $signed(hiddenLayer_43) * $signed(io_weightVec_43); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1844 = $signed(hiddenLayer_44) * $signed(io_weightVec_44); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1845 = $signed(hiddenLayer_45) * $signed(io_weightVec_45); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1846 = $signed(hiddenLayer_46) * $signed(io_weightVec_46); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1847 = $signed(hiddenLayer_47) * $signed(io_weightVec_47); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1848 = $signed(hiddenLayer_48) * $signed(io_weightVec_48); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1849 = $signed(hiddenLayer_49) * $signed(io_weightVec_49); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1850 = $signed(hiddenLayer_50) * $signed(io_weightVec_50); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1851 = $signed(hiddenLayer_51) * $signed(io_weightVec_51); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1852 = $signed(hiddenLayer_52) * $signed(io_weightVec_52); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1853 = $signed(hiddenLayer_53) * $signed(io_weightVec_53); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1854 = $signed(hiddenLayer_54) * $signed(io_weightVec_54); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1855 = $signed(hiddenLayer_55) * $signed(io_weightVec_55); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1856 = $signed(hiddenLayer_56) * $signed(io_weightVec_56); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1857 = $signed(hiddenLayer_57) * $signed(io_weightVec_57); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1858 = $signed(hiddenLayer_58) * $signed(io_weightVec_58); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1859 = $signed(hiddenLayer_59) * $signed(io_weightVec_59); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1860 = $signed(hiddenLayer_60) * $signed(io_weightVec_60); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1861 = $signed(hiddenLayer_61) * $signed(io_weightVec_61); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1862 = $signed(hiddenLayer_62) * $signed(io_weightVec_62); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1863 = $signed(hiddenLayer_63) * $signed(io_weightVec_63); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1864 = $signed(hiddenLayer_64) * $signed(io_weightVec_64); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1865 = $signed(hiddenLayer_65) * $signed(io_weightVec_65); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1866 = $signed(hiddenLayer_66) * $signed(io_weightVec_66); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1867 = $signed(hiddenLayer_67) * $signed(io_weightVec_67); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1868 = $signed(hiddenLayer_68) * $signed(io_weightVec_68); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1869 = $signed(hiddenLayer_69) * $signed(io_weightVec_69); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1870 = $signed(hiddenLayer_70) * $signed(io_weightVec_70); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1871 = $signed(hiddenLayer_71) * $signed(io_weightVec_71); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1872 = $signed(hiddenLayer_72) * $signed(io_weightVec_72); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1873 = $signed(hiddenLayer_73) * $signed(io_weightVec_73); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1874 = $signed(hiddenLayer_74) * $signed(io_weightVec_74); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1875 = $signed(hiddenLayer_75) * $signed(io_weightVec_75); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1876 = $signed(hiddenLayer_76) * $signed(io_weightVec_76); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1877 = $signed(hiddenLayer_77) * $signed(io_weightVec_77); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1878 = $signed(hiddenLayer_78) * $signed(io_weightVec_78); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1879 = $signed(hiddenLayer_79) * $signed(io_weightVec_79); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1880 = $signed(hiddenLayer_80) * $signed(io_weightVec_80); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1881 = $signed(hiddenLayer_81) * $signed(io_weightVec_81); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1882 = $signed(hiddenLayer_82) * $signed(io_weightVec_82); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1883 = $signed(hiddenLayer_83) * $signed(io_weightVec_83); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1884 = $signed(hiddenLayer_84) * $signed(io_weightVec_84); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1885 = $signed(hiddenLayer_85) * $signed(io_weightVec_85); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1886 = $signed(hiddenLayer_86) * $signed(io_weightVec_86); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1887 = $signed(hiddenLayer_87) * $signed(io_weightVec_87); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1888 = $signed(hiddenLayer_88) * $signed(io_weightVec_88); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1889 = $signed(hiddenLayer_89) * $signed(io_weightVec_89); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1890 = $signed(hiddenLayer_90) * $signed(io_weightVec_90); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1891 = $signed(hiddenLayer_91) * $signed(io_weightVec_91); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1892 = $signed(hiddenLayer_92) * $signed(io_weightVec_92); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1893 = $signed(hiddenLayer_93) * $signed(io_weightVec_93); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1894 = $signed(hiddenLayer_94) * $signed(io_weightVec_94); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1895 = $signed(hiddenLayer_95) * $signed(io_weightVec_95); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1896 = $signed(hiddenLayer_96) * $signed(io_weightVec_96); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1897 = $signed(hiddenLayer_97) * $signed(io_weightVec_97); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1898 = $signed(hiddenLayer_98) * $signed(io_weightVec_98); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1899 = $signed(hiddenLayer_99) * $signed(io_weightVec_99); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1901 = $signed(_T_1800) + $signed(_T_1801); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1902 = $signed(_T_1901); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1904 = $signed(_T_1902) + $signed(_T_1802); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1905 = $signed(_T_1904); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1907 = $signed(_T_1905) + $signed(_T_1803); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1908 = $signed(_T_1907); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1910 = $signed(_T_1908) + $signed(_T_1804); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1911 = $signed(_T_1910); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1913 = $signed(_T_1911) + $signed(_T_1805); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1914 = $signed(_T_1913); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1916 = $signed(_T_1914) + $signed(_T_1806); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1917 = $signed(_T_1916); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1919 = $signed(_T_1917) + $signed(_T_1807); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1920 = $signed(_T_1919); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1922 = $signed(_T_1920) + $signed(_T_1808); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1923 = $signed(_T_1922); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1925 = $signed(_T_1923) + $signed(_T_1809); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1926 = $signed(_T_1925); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1928 = $signed(_T_1926) + $signed(_T_1810); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1929 = $signed(_T_1928); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1931 = $signed(_T_1929) + $signed(_T_1811); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1932 = $signed(_T_1931); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1934 = $signed(_T_1932) + $signed(_T_1812); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1935 = $signed(_T_1934); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1937 = $signed(_T_1935) + $signed(_T_1813); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1938 = $signed(_T_1937); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1940 = $signed(_T_1938) + $signed(_T_1814); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1941 = $signed(_T_1940); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1943 = $signed(_T_1941) + $signed(_T_1815); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1944 = $signed(_T_1943); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1946 = $signed(_T_1944) + $signed(_T_1816); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1947 = $signed(_T_1946); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1949 = $signed(_T_1947) + $signed(_T_1817); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1950 = $signed(_T_1949); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1952 = $signed(_T_1950) + $signed(_T_1818); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1953 = $signed(_T_1952); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1955 = $signed(_T_1953) + $signed(_T_1819); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1956 = $signed(_T_1955); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1958 = $signed(_T_1956) + $signed(_T_1820); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1959 = $signed(_T_1958); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1961 = $signed(_T_1959) + $signed(_T_1821); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1962 = $signed(_T_1961); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1964 = $signed(_T_1962) + $signed(_T_1822); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1965 = $signed(_T_1964); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1967 = $signed(_T_1965) + $signed(_T_1823); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1968 = $signed(_T_1967); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1970 = $signed(_T_1968) + $signed(_T_1824); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1971 = $signed(_T_1970); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1973 = $signed(_T_1971) + $signed(_T_1825); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1974 = $signed(_T_1973); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1976 = $signed(_T_1974) + $signed(_T_1826); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1977 = $signed(_T_1976); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1979 = $signed(_T_1977) + $signed(_T_1827); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1980 = $signed(_T_1979); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1982 = $signed(_T_1980) + $signed(_T_1828); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1983 = $signed(_T_1982); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1985 = $signed(_T_1983) + $signed(_T_1829); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1986 = $signed(_T_1985); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1988 = $signed(_T_1986) + $signed(_T_1830); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1989 = $signed(_T_1988); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1991 = $signed(_T_1989) + $signed(_T_1831); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1992 = $signed(_T_1991); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1994 = $signed(_T_1992) + $signed(_T_1832); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1995 = $signed(_T_1994); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1997 = $signed(_T_1995) + $signed(_T_1833); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1998 = $signed(_T_1997); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2000 = $signed(_T_1998) + $signed(_T_1834); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2001 = $signed(_T_2000); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2003 = $signed(_T_2001) + $signed(_T_1835); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2004 = $signed(_T_2003); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2006 = $signed(_T_2004) + $signed(_T_1836); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2007 = $signed(_T_2006); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2009 = $signed(_T_2007) + $signed(_T_1837); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2010 = $signed(_T_2009); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2012 = $signed(_T_2010) + $signed(_T_1838); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2013 = $signed(_T_2012); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2015 = $signed(_T_2013) + $signed(_T_1839); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2016 = $signed(_T_2015); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2018 = $signed(_T_2016) + $signed(_T_1840); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2019 = $signed(_T_2018); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2021 = $signed(_T_2019) + $signed(_T_1841); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2022 = $signed(_T_2021); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2024 = $signed(_T_2022) + $signed(_T_1842); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2025 = $signed(_T_2024); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2027 = $signed(_T_2025) + $signed(_T_1843); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2028 = $signed(_T_2027); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2030 = $signed(_T_2028) + $signed(_T_1844); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2031 = $signed(_T_2030); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2033 = $signed(_T_2031) + $signed(_T_1845); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2034 = $signed(_T_2033); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2036 = $signed(_T_2034) + $signed(_T_1846); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2037 = $signed(_T_2036); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2039 = $signed(_T_2037) + $signed(_T_1847); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2040 = $signed(_T_2039); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2042 = $signed(_T_2040) + $signed(_T_1848); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2043 = $signed(_T_2042); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2045 = $signed(_T_2043) + $signed(_T_1849); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2046 = $signed(_T_2045); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2048 = $signed(_T_2046) + $signed(_T_1850); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2049 = $signed(_T_2048); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2051 = $signed(_T_2049) + $signed(_T_1851); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2052 = $signed(_T_2051); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2054 = $signed(_T_2052) + $signed(_T_1852); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2055 = $signed(_T_2054); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2057 = $signed(_T_2055) + $signed(_T_1853); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2058 = $signed(_T_2057); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2060 = $signed(_T_2058) + $signed(_T_1854); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2061 = $signed(_T_2060); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2063 = $signed(_T_2061) + $signed(_T_1855); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2064 = $signed(_T_2063); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2066 = $signed(_T_2064) + $signed(_T_1856); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2067 = $signed(_T_2066); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2069 = $signed(_T_2067) + $signed(_T_1857); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2070 = $signed(_T_2069); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2072 = $signed(_T_2070) + $signed(_T_1858); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2073 = $signed(_T_2072); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2075 = $signed(_T_2073) + $signed(_T_1859); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2076 = $signed(_T_2075); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2078 = $signed(_T_2076) + $signed(_T_1860); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2079 = $signed(_T_2078); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2081 = $signed(_T_2079) + $signed(_T_1861); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2082 = $signed(_T_2081); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2084 = $signed(_T_2082) + $signed(_T_1862); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2085 = $signed(_T_2084); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2087 = $signed(_T_2085) + $signed(_T_1863); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2088 = $signed(_T_2087); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2090 = $signed(_T_2088) + $signed(_T_1864); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2091 = $signed(_T_2090); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2093 = $signed(_T_2091) + $signed(_T_1865); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2094 = $signed(_T_2093); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2096 = $signed(_T_2094) + $signed(_T_1866); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2097 = $signed(_T_2096); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2099 = $signed(_T_2097) + $signed(_T_1867); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2100 = $signed(_T_2099); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2102 = $signed(_T_2100) + $signed(_T_1868); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2103 = $signed(_T_2102); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2105 = $signed(_T_2103) + $signed(_T_1869); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2106 = $signed(_T_2105); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2108 = $signed(_T_2106) + $signed(_T_1870); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2109 = $signed(_T_2108); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2111 = $signed(_T_2109) + $signed(_T_1871); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2112 = $signed(_T_2111); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2114 = $signed(_T_2112) + $signed(_T_1872); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2115 = $signed(_T_2114); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2117 = $signed(_T_2115) + $signed(_T_1873); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2118 = $signed(_T_2117); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2120 = $signed(_T_2118) + $signed(_T_1874); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2121 = $signed(_T_2120); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2123 = $signed(_T_2121) + $signed(_T_1875); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2124 = $signed(_T_2123); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2126 = $signed(_T_2124) + $signed(_T_1876); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2127 = $signed(_T_2126); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2129 = $signed(_T_2127) + $signed(_T_1877); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2130 = $signed(_T_2129); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2132 = $signed(_T_2130) + $signed(_T_1878); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2133 = $signed(_T_2132); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2135 = $signed(_T_2133) + $signed(_T_1879); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2136 = $signed(_T_2135); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2138 = $signed(_T_2136) + $signed(_T_1880); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2139 = $signed(_T_2138); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2141 = $signed(_T_2139) + $signed(_T_1881); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2142 = $signed(_T_2141); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2144 = $signed(_T_2142) + $signed(_T_1882); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2145 = $signed(_T_2144); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2147 = $signed(_T_2145) + $signed(_T_1883); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2148 = $signed(_T_2147); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2150 = $signed(_T_2148) + $signed(_T_1884); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2151 = $signed(_T_2150); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2153 = $signed(_T_2151) + $signed(_T_1885); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2154 = $signed(_T_2153); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2156 = $signed(_T_2154) + $signed(_T_1886); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2157 = $signed(_T_2156); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2159 = $signed(_T_2157) + $signed(_T_1887); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2160 = $signed(_T_2159); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2162 = $signed(_T_2160) + $signed(_T_1888); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2163 = $signed(_T_2162); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2165 = $signed(_T_2163) + $signed(_T_1889); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2166 = $signed(_T_2165); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2168 = $signed(_T_2166) + $signed(_T_1890); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2169 = $signed(_T_2168); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2171 = $signed(_T_2169) + $signed(_T_1891); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2172 = $signed(_T_2171); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2174 = $signed(_T_2172) + $signed(_T_1892); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2175 = $signed(_T_2174); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2177 = $signed(_T_2175) + $signed(_T_1893); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2178 = $signed(_T_2177); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2180 = $signed(_T_2178) + $signed(_T_1894); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2181 = $signed(_T_2180); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2183 = $signed(_T_2181) + $signed(_T_1895); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2184 = $signed(_T_2183); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2186 = $signed(_T_2184) + $signed(_T_1896); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2187 = $signed(_T_2186); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2189 = $signed(_T_2187) + $signed(_T_1897); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2190 = $signed(_T_2189); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2192 = $signed(_T_2190) + $signed(_T_1898); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2193 = $signed(_T_2192); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2195 = $signed(_T_2193) + $signed(_T_1899); // @[FixedPointTypeClass.scala 21:58]
  assign _T_2196 = $signed(_T_2195); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_202 = _T_2196[63:8]; // @[neuralNet.scala 66:24 neuralNet.scala 68:16 neuralNet.scala 68:16 neuralNet.scala 68:16 neuralNet.scala 68:16]
  assign _GEN_203 = _GEN_202[31:0]; // @[neuralNet.scala 66:24 neuralNet.scala 68:16 neuralNet.scala 68:16 neuralNet.scala 68:16 neuralNet.scala 68:16]
  assign dotProduct = $signed(_GEN_203); // @[neuralNet.scala 66:24 neuralNet.scala 68:16 neuralNet.scala 68:16 neuralNet.scala 68:16 neuralNet.scala 68:16]
  assign _T_3389 = $signed(dotProduct) + $signed(io_biasScalar); // @[FixedPointTypeClass.scala 21:58]
  assign actualPreReLU = $signed(_T_3389); // @[FixedPointTypeClass.scala 21:58]
  assign _T_3391 = $signed(actualPreReLU) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign actualVotes = _T_3391 ? $signed(actualPreReLU) : $signed(32'sh0); // @[neuralNet.scala 75:21]
  assign finalPredict = $signed(actualVotes) > $signed(32'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign io_out_valid = valReg; // @[neuralNet.scala 89:16]
  assign io_out_bits = outReg; // @[neuralNet.scala 88:15]
  assign io_rawVotes = rawVotesReg; // @[neuralNet.scala 87:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  rawVotesReg = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  outReg = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  valReg = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (io_in_valid) begin
      if (_T_3391) begin
        rawVotesReg <= actualPreReLU;
      end else begin
        rawVotesReg <= 32'sh0;
      end
    end
    if (io_in_valid) begin
      outReg <= finalPredict;
    end
    valReg <= io_in_valid;
  end
endmodule
module WellnessModule(
  input         clock,
  input         reset,
  input         io_streamIn_valid,
  input  [31:0] io_streamIn_bits,
  input         io_in_valid,
  input  [31:0] io_in_bits,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_0_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_0_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_0_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_0_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_1_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_1_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_1_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_1_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_2_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_2_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_2_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_2_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_3_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_3_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_3_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_3_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_4_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_4_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_4_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_4_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_5_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_5_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_5_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_5_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_6_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_6_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_6_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_6_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_7_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_7_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_7_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_7_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_8_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_8_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_8_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_8_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_9_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_9_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_9_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_9_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_10_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_10_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_10_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_10_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_11_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_11_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_11_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_11_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_12_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_12_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_12_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_12_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_13_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_13_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_13_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_13_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_14_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_14_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_14_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_14_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_15_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_15_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_15_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_15_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_16_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_16_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_16_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_16_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_17_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_17_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_17_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_17_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_18_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_18_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_18_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_18_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_19_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_19_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_19_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_19_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_20_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_20_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_20_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_20_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_21_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_21_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_21_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_21_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_22_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_22_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_22_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_22_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_23_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_23_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_23_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_23_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_24_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_24_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_24_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_24_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_25_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_25_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_25_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_25_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_26_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_26_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_26_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_26_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_27_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_27_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_27_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_27_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_28_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_28_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_28_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_28_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_29_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_29_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_29_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_29_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_30_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_30_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_30_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_30_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_31_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_31_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_31_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_31_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_32_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_32_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_32_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_32_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_33_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_33_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_33_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_33_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_34_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_34_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_34_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_34_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_35_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_35_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_35_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_35_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_36_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_36_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_36_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_36_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_37_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_37_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_37_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_37_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_38_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_38_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_38_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_38_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_39_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_39_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_39_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_39_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_40_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_40_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_40_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_40_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_41_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_41_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_41_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_41_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_42_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_42_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_42_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_42_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_43_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_43_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_43_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_43_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_44_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_44_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_44_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_44_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_45_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_45_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_45_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_45_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_46_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_46_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_46_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_46_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_47_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_47_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_47_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_47_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_48_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_48_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_48_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_48_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_49_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_49_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_49_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_49_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_50_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_50_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_50_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_50_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_51_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_51_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_51_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_51_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_52_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_52_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_52_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_52_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_53_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_53_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_53_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_53_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_54_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_54_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_54_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_54_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_55_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_55_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_55_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_55_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_56_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_56_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_56_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_56_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_57_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_57_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_57_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_57_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_58_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_58_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_58_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_58_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_59_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_59_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_59_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_59_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_60_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_60_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_60_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_60_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_61_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_61_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_61_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_61_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_62_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_62_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_62_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_62_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_63_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_63_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_63_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_63_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_64_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_64_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_64_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_64_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_65_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_65_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_65_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_65_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_66_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_66_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_66_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_66_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_67_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_67_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_67_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_67_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_68_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_68_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_68_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_68_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_69_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_69_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_69_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_69_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_70_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_70_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_70_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_70_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_71_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_71_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_71_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_71_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_72_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_72_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_72_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_72_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_73_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_73_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_73_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_73_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_74_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_74_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_74_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_74_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_75_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_75_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_75_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_75_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_76_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_76_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_76_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_76_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_77_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_77_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_77_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_77_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_78_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_78_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_78_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_78_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_79_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_79_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_79_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_79_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_80_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_80_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_80_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_80_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_81_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_81_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_81_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_81_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_82_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_82_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_82_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_82_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_83_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_83_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_83_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_83_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_84_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_84_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_84_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_84_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_85_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_85_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_85_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_85_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_86_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_86_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_86_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_86_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_87_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_87_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_87_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_87_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_88_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_88_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_88_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_88_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_89_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_89_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_89_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_89_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_90_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_90_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_90_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_90_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_91_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_91_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_91_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_91_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_92_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_92_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_92_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_92_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_93_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_93_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_93_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_93_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_94_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_94_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_94_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_94_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_95_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_95_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_95_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_95_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_96_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_96_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_96_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_96_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_97_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_97_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_97_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_97_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_98_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_98_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_98_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_98_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_99_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_99_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_99_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightMatrix_99_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_0,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_1,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_2,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_3,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_4,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_5,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_6,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_7,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_8,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_9,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_10,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_11,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_12,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_13,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_14,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_15,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_16,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_17,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_18,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_19,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_20,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_21,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_22,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_23,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_24,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_25,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_26,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_27,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_28,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_29,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_30,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_31,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_32,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_33,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_34,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_35,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_36,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_37,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_38,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_39,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_40,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_41,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_42,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_43,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_44,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_45,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_46,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_47,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_48,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_49,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_50,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_51,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_52,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_53,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_54,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_55,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_56,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_57,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_58,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_59,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_60,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_61,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_62,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_63,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_64,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_65,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_66,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_67,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_68,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_69,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_70,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_71,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_72,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_73,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_74,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_75,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_76,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_77,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_78,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_79,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_80,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_81,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_82,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_83,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_84,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_85,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_86,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_87,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_88,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_89,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_90,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_91,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_92,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_93,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_94,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_95,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_96,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_97,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_98,
  input  [31:0] io_inConf_bits_confneuralNetsweightVec_99,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_0,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_1,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_2,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_3,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_4,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_5,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_6,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_7,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_8,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_9,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_10,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_11,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_12,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_13,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_14,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_15,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_16,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_17,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_18,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_19,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_20,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_21,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_22,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_23,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_24,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_25,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_26,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_27,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_28,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_29,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_30,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_31,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_32,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_33,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_34,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_35,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_36,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_37,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_38,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_39,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_40,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_41,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_42,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_43,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_44,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_45,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_46,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_47,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_48,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_49,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_50,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_51,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_52,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_53,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_54,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_55,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_56,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_57,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_58,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_59,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_60,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_61,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_62,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_63,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_64,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_65,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_66,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_67,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_68,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_69,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_70,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_71,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_72,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_73,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_74,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_75,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_76,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_77,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_78,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_79,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_80,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_81,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_82,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_83,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_84,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_85,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_86,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_87,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_88,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_89,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_90,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_91,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_92,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_93,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_94,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_95,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_96,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_97,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_98,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVec_99,
  input  [31:0] io_inConf_bits_confneuralNetsbiasScalar_0,
  input         io_inConf_bits_confInputMuxSel,
  output        io_out_valid,
  output        io_out_bits,
  output [31:0] io_rawVotes
);
  wire  filter1_clock; // @[Wellness.scala 255:23]
  wire  filter1_reset; // @[Wellness.scala 255:23]
  wire  filter1_io_in_valid; // @[Wellness.scala 255:23]
  wire [31:0] filter1_io_in_bits; // @[Wellness.scala 255:23]
  wire  filter1_io_out_valid; // @[Wellness.scala 255:23]
  wire [31:0] filter1_io_out_bits; // @[Wellness.scala 255:23]
  wire  lineLength1_clock; // @[Wellness.scala 256:27]
  wire  lineLength1_reset; // @[Wellness.scala 256:27]
  wire  lineLength1_io_in_valid; // @[Wellness.scala 256:27]
  wire [31:0] lineLength1_io_in_bits; // @[Wellness.scala 256:27]
  wire  lineLength1_io_out_valid; // @[Wellness.scala 256:27]
  wire [31:0] lineLength1_io_out_bits; // @[Wellness.scala 256:27]
  wire  filterAlpha_clock; // @[Wellness.scala 258:27]
  wire  filterAlpha_reset; // @[Wellness.scala 258:27]
  wire  filterAlpha_io_in_valid; // @[Wellness.scala 258:27]
  wire [31:0] filterAlpha_io_in_bits; // @[Wellness.scala 258:27]
  wire  filterAlpha_io_out_valid; // @[Wellness.scala 258:27]
  wire [31:0] filterAlpha_io_out_bits; // @[Wellness.scala 258:27]
  wire  filterBeta_clock; // @[Wellness.scala 259:26]
  wire  filterBeta_reset; // @[Wellness.scala 259:26]
  wire  filterBeta_io_in_valid; // @[Wellness.scala 259:26]
  wire [31:0] filterBeta_io_in_bits; // @[Wellness.scala 259:26]
  wire  filterBeta_io_out_valid; // @[Wellness.scala 259:26]
  wire [31:0] filterBeta_io_out_bits; // @[Wellness.scala 259:26]
  wire  filterGamma_clock; // @[Wellness.scala 260:27]
  wire  filterGamma_reset; // @[Wellness.scala 260:27]
  wire  filterGamma_io_in_valid; // @[Wellness.scala 260:27]
  wire [31:0] filterGamma_io_in_bits; // @[Wellness.scala 260:27]
  wire  filterGamma_io_out_valid; // @[Wellness.scala 260:27]
  wire [31:0] filterGamma_io_out_bits; // @[Wellness.scala 260:27]
  wire  bandpowerAlpha_clock; // @[Wellness.scala 262:30]
  wire  bandpowerAlpha_reset; // @[Wellness.scala 262:30]
  wire  bandpowerAlpha_io_in_valid; // @[Wellness.scala 262:30]
  wire [31:0] bandpowerAlpha_io_in_bits; // @[Wellness.scala 262:30]
  wire  bandpowerAlpha_io_out_valid; // @[Wellness.scala 262:30]
  wire [31:0] bandpowerAlpha_io_out_bits; // @[Wellness.scala 262:30]
  wire  bandpowerBeta_clock; // @[Wellness.scala 263:29]
  wire  bandpowerBeta_reset; // @[Wellness.scala 263:29]
  wire  bandpowerBeta_io_in_valid; // @[Wellness.scala 263:29]
  wire [31:0] bandpowerBeta_io_in_bits; // @[Wellness.scala 263:29]
  wire  bandpowerBeta_io_out_valid; // @[Wellness.scala 263:29]
  wire [31:0] bandpowerBeta_io_out_bits; // @[Wellness.scala 263:29]
  wire  bandpowerGamma_clock; // @[Wellness.scala 264:30]
  wire  bandpowerGamma_reset; // @[Wellness.scala 264:30]
  wire  bandpowerGamma_io_in_valid; // @[Wellness.scala 264:30]
  wire [31:0] bandpowerGamma_io_in_bits; // @[Wellness.scala 264:30]
  wire  bandpowerGamma_io_out_valid; // @[Wellness.scala 264:30]
  wire [31:0] bandpowerGamma_io_out_bits; // @[Wellness.scala 264:30]
  wire  neuralNets_clock; // @[Wellness.scala 266:26]
  wire  neuralNets_io_in_valid; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_in_bits_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_in_bits_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_in_bits_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_in_bits_3; // @[Wellness.scala 266:26]
  wire  neuralNets_io_out_valid; // @[Wellness.scala 266:26]
  wire  neuralNets_io_out_bits; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_0_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_0_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_0_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_0_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_1_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_1_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_1_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_1_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_2_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_2_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_2_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_2_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_3_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_3_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_3_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_3_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_4_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_4_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_4_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_4_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_5_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_5_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_5_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_5_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_6_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_6_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_6_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_6_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_7_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_7_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_7_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_7_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_8_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_8_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_8_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_8_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_9_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_9_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_9_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_9_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_10_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_10_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_10_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_10_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_11_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_11_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_11_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_11_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_12_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_12_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_12_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_12_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_13_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_13_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_13_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_13_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_14_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_14_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_14_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_14_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_15_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_15_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_15_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_15_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_16_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_16_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_16_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_16_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_17_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_17_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_17_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_17_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_18_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_18_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_18_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_18_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_19_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_19_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_19_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_19_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_20_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_20_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_20_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_20_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_21_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_21_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_21_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_21_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_22_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_22_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_22_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_22_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_23_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_23_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_23_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_23_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_24_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_24_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_24_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_24_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_25_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_25_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_25_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_25_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_26_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_26_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_26_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_26_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_27_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_27_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_27_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_27_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_28_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_28_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_28_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_28_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_29_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_29_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_29_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_29_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_30_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_30_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_30_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_30_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_31_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_31_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_31_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_31_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_32_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_32_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_32_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_32_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_33_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_33_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_33_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_33_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_34_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_34_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_34_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_34_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_35_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_35_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_35_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_35_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_36_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_36_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_36_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_36_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_37_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_37_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_37_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_37_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_38_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_38_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_38_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_38_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_39_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_39_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_39_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_39_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_40_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_40_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_40_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_40_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_41_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_41_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_41_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_41_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_42_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_42_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_42_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_42_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_43_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_43_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_43_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_43_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_44_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_44_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_44_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_44_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_45_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_45_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_45_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_45_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_46_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_46_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_46_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_46_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_47_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_47_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_47_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_47_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_48_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_48_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_48_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_48_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_49_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_49_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_49_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_49_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_50_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_50_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_50_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_50_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_51_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_51_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_51_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_51_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_52_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_52_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_52_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_52_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_53_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_53_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_53_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_53_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_54_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_54_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_54_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_54_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_55_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_55_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_55_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_55_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_56_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_56_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_56_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_56_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_57_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_57_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_57_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_57_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_58_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_58_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_58_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_58_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_59_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_59_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_59_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_59_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_60_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_60_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_60_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_60_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_61_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_61_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_61_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_61_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_62_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_62_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_62_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_62_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_63_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_63_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_63_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_63_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_64_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_64_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_64_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_64_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_65_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_65_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_65_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_65_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_66_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_66_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_66_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_66_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_67_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_67_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_67_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_67_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_68_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_68_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_68_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_68_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_69_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_69_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_69_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_69_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_70_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_70_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_70_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_70_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_71_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_71_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_71_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_71_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_72_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_72_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_72_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_72_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_73_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_73_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_73_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_73_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_74_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_74_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_74_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_74_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_75_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_75_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_75_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_75_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_76_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_76_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_76_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_76_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_77_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_77_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_77_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_77_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_78_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_78_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_78_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_78_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_79_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_79_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_79_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_79_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_80_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_80_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_80_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_80_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_81_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_81_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_81_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_81_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_82_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_82_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_82_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_82_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_83_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_83_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_83_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_83_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_84_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_84_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_84_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_84_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_85_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_85_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_85_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_85_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_86_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_86_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_86_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_86_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_87_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_87_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_87_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_87_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_88_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_88_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_88_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_88_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_89_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_89_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_89_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_89_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_90_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_90_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_90_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_90_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_91_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_91_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_91_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_91_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_92_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_92_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_92_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_92_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_93_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_93_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_93_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_93_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_94_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_94_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_94_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_94_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_95_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_95_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_95_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_95_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_96_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_96_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_96_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_96_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_97_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_97_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_97_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_97_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_98_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_98_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_98_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_98_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_99_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_99_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_99_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightMatrix_99_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_4; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_5; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_6; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_7; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_8; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_9; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_10; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_11; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_12; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_13; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_14; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_15; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_16; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_17; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_18; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_19; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_20; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_21; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_22; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_23; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_24; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_25; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_26; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_27; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_28; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_29; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_30; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_31; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_32; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_33; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_34; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_35; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_36; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_37; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_38; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_39; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_40; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_41; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_42; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_43; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_44; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_45; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_46; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_47; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_48; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_49; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_50; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_51; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_52; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_53; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_54; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_55; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_56; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_57; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_58; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_59; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_60; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_61; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_62; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_63; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_64; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_65; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_66; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_67; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_68; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_69; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_70; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_71; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_72; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_73; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_74; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_75; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_76; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_77; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_78; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_79; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_80; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_81; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_82; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_83; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_84; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_85; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_86; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_87; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_88; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_89; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_90; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_91; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_92; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_93; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_94; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_95; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_96; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_97; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_98; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_weightVec_99; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_4; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_5; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_6; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_7; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_8; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_9; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_10; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_11; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_12; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_13; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_14; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_15; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_16; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_17; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_18; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_19; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_20; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_21; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_22; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_23; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_24; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_25; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_26; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_27; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_28; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_29; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_30; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_31; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_32; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_33; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_34; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_35; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_36; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_37; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_38; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_39; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_40; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_41; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_42; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_43; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_44; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_45; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_46; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_47; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_48; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_49; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_50; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_51; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_52; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_53; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_54; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_55; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_56; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_57; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_58; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_59; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_60; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_61; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_62; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_63; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_64; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_65; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_66; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_67; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_68; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_69; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_70; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_71; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_72; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_73; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_74; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_75; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_76; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_77; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_78; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_79; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_80; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_81; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_82; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_83; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_84; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_85; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_86; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_87; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_88; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_89; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_90; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_91; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_92; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_93; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_94; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_95; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_96; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_97; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_98; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVec_99; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasScalar; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_rawVotes; // @[Wellness.scala 266:26]
  wire [31:0] _T_1; // @[Wellness.scala 271:80]
  wire [31:0] _T_2; // @[Wellness.scala 271:80]
  wire [31:0] _T_4; // @[Wellness.scala 271:125]
  wire [31:0] _T_5; // @[Wellness.scala 271:125]
  wire [31:0] _T_10; // @[Wellness.scala 283:57]
  wire [31:0] _T_22; // @[Wellness.scala 314:65]
  reg [31:0] lineLength1Reg1; // @[Wellness.scala 314:32]
  reg [31:0] _RAND_0;
  reg  lineLength1Valid1; // @[Wellness.scala 316:34]
  reg [31:0] _RAND_1;
  wire [31:0] _T_25; // @[Wellness.scala 327:58]
  wire [31:0] _T_28; // @[Wellness.scala 328:57]
  wire [31:0] _T_31; // @[Wellness.scala 329:58]
  wire [31:0] _T_34; // @[Wellness.scala 330:47]
  wire  _T_36; // @[Wellness.scala 332:48]
  wire  _T_37; // @[Wellness.scala 332:79]
  ConstantCoefficientFIRFilter filter1 ( // @[Wellness.scala 255:23]
    .clock(filter1_clock),
    .reset(filter1_reset),
    .io_in_valid(filter1_io_in_valid),
    .io_in_bits(filter1_io_in_bits),
    .io_out_valid(filter1_io_out_valid),
    .io_out_bits(filter1_io_out_bits)
  );
  lineLength lineLength1 ( // @[Wellness.scala 256:27]
    .clock(lineLength1_clock),
    .reset(lineLength1_reset),
    .io_in_valid(lineLength1_io_in_valid),
    .io_in_bits(lineLength1_io_in_bits),
    .io_out_valid(lineLength1_io_out_valid),
    .io_out_bits(lineLength1_io_out_bits)
  );
  ConstantCoefficientFIRFilter filterAlpha ( // @[Wellness.scala 258:27]
    .clock(filterAlpha_clock),
    .reset(filterAlpha_reset),
    .io_in_valid(filterAlpha_io_in_valid),
    .io_in_bits(filterAlpha_io_in_bits),
    .io_out_valid(filterAlpha_io_out_valid),
    .io_out_bits(filterAlpha_io_out_bits)
  );
  ConstantCoefficientFIRFilter filterBeta ( // @[Wellness.scala 259:26]
    .clock(filterBeta_clock),
    .reset(filterBeta_reset),
    .io_in_valid(filterBeta_io_in_valid),
    .io_in_bits(filterBeta_io_in_bits),
    .io_out_valid(filterBeta_io_out_valid),
    .io_out_bits(filterBeta_io_out_bits)
  );
  ConstantCoefficientFIRFilter filterGamma ( // @[Wellness.scala 260:27]
    .clock(filterGamma_clock),
    .reset(filterGamma_reset),
    .io_in_valid(filterGamma_io_in_valid),
    .io_in_bits(filterGamma_io_in_bits),
    .io_out_valid(filterGamma_io_out_valid),
    .io_out_bits(filterGamma_io_out_bits)
  );
  sumSquares bandpowerAlpha ( // @[Wellness.scala 262:30]
    .clock(bandpowerAlpha_clock),
    .reset(bandpowerAlpha_reset),
    .io_in_valid(bandpowerAlpha_io_in_valid),
    .io_in_bits(bandpowerAlpha_io_in_bits),
    .io_out_valid(bandpowerAlpha_io_out_valid),
    .io_out_bits(bandpowerAlpha_io_out_bits)
  );
  sumSquares bandpowerBeta ( // @[Wellness.scala 263:29]
    .clock(bandpowerBeta_clock),
    .reset(bandpowerBeta_reset),
    .io_in_valid(bandpowerBeta_io_in_valid),
    .io_in_bits(bandpowerBeta_io_in_bits),
    .io_out_valid(bandpowerBeta_io_out_valid),
    .io_out_bits(bandpowerBeta_io_out_bits)
  );
  sumSquares bandpowerGamma ( // @[Wellness.scala 264:30]
    .clock(bandpowerGamma_clock),
    .reset(bandpowerGamma_reset),
    .io_in_valid(bandpowerGamma_io_in_valid),
    .io_in_bits(bandpowerGamma_io_in_bits),
    .io_out_valid(bandpowerGamma_io_out_valid),
    .io_out_bits(bandpowerGamma_io_out_bits)
  );
  NeuralNet neuralNets ( // @[Wellness.scala 266:26]
    .clock(neuralNets_clock),
    .io_in_valid(neuralNets_io_in_valid),
    .io_in_bits_0(neuralNets_io_in_bits_0),
    .io_in_bits_1(neuralNets_io_in_bits_1),
    .io_in_bits_2(neuralNets_io_in_bits_2),
    .io_in_bits_3(neuralNets_io_in_bits_3),
    .io_out_valid(neuralNets_io_out_valid),
    .io_out_bits(neuralNets_io_out_bits),
    .io_weightMatrix_0_0(neuralNets_io_weightMatrix_0_0),
    .io_weightMatrix_0_1(neuralNets_io_weightMatrix_0_1),
    .io_weightMatrix_0_2(neuralNets_io_weightMatrix_0_2),
    .io_weightMatrix_0_3(neuralNets_io_weightMatrix_0_3),
    .io_weightMatrix_1_0(neuralNets_io_weightMatrix_1_0),
    .io_weightMatrix_1_1(neuralNets_io_weightMatrix_1_1),
    .io_weightMatrix_1_2(neuralNets_io_weightMatrix_1_2),
    .io_weightMatrix_1_3(neuralNets_io_weightMatrix_1_3),
    .io_weightMatrix_2_0(neuralNets_io_weightMatrix_2_0),
    .io_weightMatrix_2_1(neuralNets_io_weightMatrix_2_1),
    .io_weightMatrix_2_2(neuralNets_io_weightMatrix_2_2),
    .io_weightMatrix_2_3(neuralNets_io_weightMatrix_2_3),
    .io_weightMatrix_3_0(neuralNets_io_weightMatrix_3_0),
    .io_weightMatrix_3_1(neuralNets_io_weightMatrix_3_1),
    .io_weightMatrix_3_2(neuralNets_io_weightMatrix_3_2),
    .io_weightMatrix_3_3(neuralNets_io_weightMatrix_3_3),
    .io_weightMatrix_4_0(neuralNets_io_weightMatrix_4_0),
    .io_weightMatrix_4_1(neuralNets_io_weightMatrix_4_1),
    .io_weightMatrix_4_2(neuralNets_io_weightMatrix_4_2),
    .io_weightMatrix_4_3(neuralNets_io_weightMatrix_4_3),
    .io_weightMatrix_5_0(neuralNets_io_weightMatrix_5_0),
    .io_weightMatrix_5_1(neuralNets_io_weightMatrix_5_1),
    .io_weightMatrix_5_2(neuralNets_io_weightMatrix_5_2),
    .io_weightMatrix_5_3(neuralNets_io_weightMatrix_5_3),
    .io_weightMatrix_6_0(neuralNets_io_weightMatrix_6_0),
    .io_weightMatrix_6_1(neuralNets_io_weightMatrix_6_1),
    .io_weightMatrix_6_2(neuralNets_io_weightMatrix_6_2),
    .io_weightMatrix_6_3(neuralNets_io_weightMatrix_6_3),
    .io_weightMatrix_7_0(neuralNets_io_weightMatrix_7_0),
    .io_weightMatrix_7_1(neuralNets_io_weightMatrix_7_1),
    .io_weightMatrix_7_2(neuralNets_io_weightMatrix_7_2),
    .io_weightMatrix_7_3(neuralNets_io_weightMatrix_7_3),
    .io_weightMatrix_8_0(neuralNets_io_weightMatrix_8_0),
    .io_weightMatrix_8_1(neuralNets_io_weightMatrix_8_1),
    .io_weightMatrix_8_2(neuralNets_io_weightMatrix_8_2),
    .io_weightMatrix_8_3(neuralNets_io_weightMatrix_8_3),
    .io_weightMatrix_9_0(neuralNets_io_weightMatrix_9_0),
    .io_weightMatrix_9_1(neuralNets_io_weightMatrix_9_1),
    .io_weightMatrix_9_2(neuralNets_io_weightMatrix_9_2),
    .io_weightMatrix_9_3(neuralNets_io_weightMatrix_9_3),
    .io_weightMatrix_10_0(neuralNets_io_weightMatrix_10_0),
    .io_weightMatrix_10_1(neuralNets_io_weightMatrix_10_1),
    .io_weightMatrix_10_2(neuralNets_io_weightMatrix_10_2),
    .io_weightMatrix_10_3(neuralNets_io_weightMatrix_10_3),
    .io_weightMatrix_11_0(neuralNets_io_weightMatrix_11_0),
    .io_weightMatrix_11_1(neuralNets_io_weightMatrix_11_1),
    .io_weightMatrix_11_2(neuralNets_io_weightMatrix_11_2),
    .io_weightMatrix_11_3(neuralNets_io_weightMatrix_11_3),
    .io_weightMatrix_12_0(neuralNets_io_weightMatrix_12_0),
    .io_weightMatrix_12_1(neuralNets_io_weightMatrix_12_1),
    .io_weightMatrix_12_2(neuralNets_io_weightMatrix_12_2),
    .io_weightMatrix_12_3(neuralNets_io_weightMatrix_12_3),
    .io_weightMatrix_13_0(neuralNets_io_weightMatrix_13_0),
    .io_weightMatrix_13_1(neuralNets_io_weightMatrix_13_1),
    .io_weightMatrix_13_2(neuralNets_io_weightMatrix_13_2),
    .io_weightMatrix_13_3(neuralNets_io_weightMatrix_13_3),
    .io_weightMatrix_14_0(neuralNets_io_weightMatrix_14_0),
    .io_weightMatrix_14_1(neuralNets_io_weightMatrix_14_1),
    .io_weightMatrix_14_2(neuralNets_io_weightMatrix_14_2),
    .io_weightMatrix_14_3(neuralNets_io_weightMatrix_14_3),
    .io_weightMatrix_15_0(neuralNets_io_weightMatrix_15_0),
    .io_weightMatrix_15_1(neuralNets_io_weightMatrix_15_1),
    .io_weightMatrix_15_2(neuralNets_io_weightMatrix_15_2),
    .io_weightMatrix_15_3(neuralNets_io_weightMatrix_15_3),
    .io_weightMatrix_16_0(neuralNets_io_weightMatrix_16_0),
    .io_weightMatrix_16_1(neuralNets_io_weightMatrix_16_1),
    .io_weightMatrix_16_2(neuralNets_io_weightMatrix_16_2),
    .io_weightMatrix_16_3(neuralNets_io_weightMatrix_16_3),
    .io_weightMatrix_17_0(neuralNets_io_weightMatrix_17_0),
    .io_weightMatrix_17_1(neuralNets_io_weightMatrix_17_1),
    .io_weightMatrix_17_2(neuralNets_io_weightMatrix_17_2),
    .io_weightMatrix_17_3(neuralNets_io_weightMatrix_17_3),
    .io_weightMatrix_18_0(neuralNets_io_weightMatrix_18_0),
    .io_weightMatrix_18_1(neuralNets_io_weightMatrix_18_1),
    .io_weightMatrix_18_2(neuralNets_io_weightMatrix_18_2),
    .io_weightMatrix_18_3(neuralNets_io_weightMatrix_18_3),
    .io_weightMatrix_19_0(neuralNets_io_weightMatrix_19_0),
    .io_weightMatrix_19_1(neuralNets_io_weightMatrix_19_1),
    .io_weightMatrix_19_2(neuralNets_io_weightMatrix_19_2),
    .io_weightMatrix_19_3(neuralNets_io_weightMatrix_19_3),
    .io_weightMatrix_20_0(neuralNets_io_weightMatrix_20_0),
    .io_weightMatrix_20_1(neuralNets_io_weightMatrix_20_1),
    .io_weightMatrix_20_2(neuralNets_io_weightMatrix_20_2),
    .io_weightMatrix_20_3(neuralNets_io_weightMatrix_20_3),
    .io_weightMatrix_21_0(neuralNets_io_weightMatrix_21_0),
    .io_weightMatrix_21_1(neuralNets_io_weightMatrix_21_1),
    .io_weightMatrix_21_2(neuralNets_io_weightMatrix_21_2),
    .io_weightMatrix_21_3(neuralNets_io_weightMatrix_21_3),
    .io_weightMatrix_22_0(neuralNets_io_weightMatrix_22_0),
    .io_weightMatrix_22_1(neuralNets_io_weightMatrix_22_1),
    .io_weightMatrix_22_2(neuralNets_io_weightMatrix_22_2),
    .io_weightMatrix_22_3(neuralNets_io_weightMatrix_22_3),
    .io_weightMatrix_23_0(neuralNets_io_weightMatrix_23_0),
    .io_weightMatrix_23_1(neuralNets_io_weightMatrix_23_1),
    .io_weightMatrix_23_2(neuralNets_io_weightMatrix_23_2),
    .io_weightMatrix_23_3(neuralNets_io_weightMatrix_23_3),
    .io_weightMatrix_24_0(neuralNets_io_weightMatrix_24_0),
    .io_weightMatrix_24_1(neuralNets_io_weightMatrix_24_1),
    .io_weightMatrix_24_2(neuralNets_io_weightMatrix_24_2),
    .io_weightMatrix_24_3(neuralNets_io_weightMatrix_24_3),
    .io_weightMatrix_25_0(neuralNets_io_weightMatrix_25_0),
    .io_weightMatrix_25_1(neuralNets_io_weightMatrix_25_1),
    .io_weightMatrix_25_2(neuralNets_io_weightMatrix_25_2),
    .io_weightMatrix_25_3(neuralNets_io_weightMatrix_25_3),
    .io_weightMatrix_26_0(neuralNets_io_weightMatrix_26_0),
    .io_weightMatrix_26_1(neuralNets_io_weightMatrix_26_1),
    .io_weightMatrix_26_2(neuralNets_io_weightMatrix_26_2),
    .io_weightMatrix_26_3(neuralNets_io_weightMatrix_26_3),
    .io_weightMatrix_27_0(neuralNets_io_weightMatrix_27_0),
    .io_weightMatrix_27_1(neuralNets_io_weightMatrix_27_1),
    .io_weightMatrix_27_2(neuralNets_io_weightMatrix_27_2),
    .io_weightMatrix_27_3(neuralNets_io_weightMatrix_27_3),
    .io_weightMatrix_28_0(neuralNets_io_weightMatrix_28_0),
    .io_weightMatrix_28_1(neuralNets_io_weightMatrix_28_1),
    .io_weightMatrix_28_2(neuralNets_io_weightMatrix_28_2),
    .io_weightMatrix_28_3(neuralNets_io_weightMatrix_28_3),
    .io_weightMatrix_29_0(neuralNets_io_weightMatrix_29_0),
    .io_weightMatrix_29_1(neuralNets_io_weightMatrix_29_1),
    .io_weightMatrix_29_2(neuralNets_io_weightMatrix_29_2),
    .io_weightMatrix_29_3(neuralNets_io_weightMatrix_29_3),
    .io_weightMatrix_30_0(neuralNets_io_weightMatrix_30_0),
    .io_weightMatrix_30_1(neuralNets_io_weightMatrix_30_1),
    .io_weightMatrix_30_2(neuralNets_io_weightMatrix_30_2),
    .io_weightMatrix_30_3(neuralNets_io_weightMatrix_30_3),
    .io_weightMatrix_31_0(neuralNets_io_weightMatrix_31_0),
    .io_weightMatrix_31_1(neuralNets_io_weightMatrix_31_1),
    .io_weightMatrix_31_2(neuralNets_io_weightMatrix_31_2),
    .io_weightMatrix_31_3(neuralNets_io_weightMatrix_31_3),
    .io_weightMatrix_32_0(neuralNets_io_weightMatrix_32_0),
    .io_weightMatrix_32_1(neuralNets_io_weightMatrix_32_1),
    .io_weightMatrix_32_2(neuralNets_io_weightMatrix_32_2),
    .io_weightMatrix_32_3(neuralNets_io_weightMatrix_32_3),
    .io_weightMatrix_33_0(neuralNets_io_weightMatrix_33_0),
    .io_weightMatrix_33_1(neuralNets_io_weightMatrix_33_1),
    .io_weightMatrix_33_2(neuralNets_io_weightMatrix_33_2),
    .io_weightMatrix_33_3(neuralNets_io_weightMatrix_33_3),
    .io_weightMatrix_34_0(neuralNets_io_weightMatrix_34_0),
    .io_weightMatrix_34_1(neuralNets_io_weightMatrix_34_1),
    .io_weightMatrix_34_2(neuralNets_io_weightMatrix_34_2),
    .io_weightMatrix_34_3(neuralNets_io_weightMatrix_34_3),
    .io_weightMatrix_35_0(neuralNets_io_weightMatrix_35_0),
    .io_weightMatrix_35_1(neuralNets_io_weightMatrix_35_1),
    .io_weightMatrix_35_2(neuralNets_io_weightMatrix_35_2),
    .io_weightMatrix_35_3(neuralNets_io_weightMatrix_35_3),
    .io_weightMatrix_36_0(neuralNets_io_weightMatrix_36_0),
    .io_weightMatrix_36_1(neuralNets_io_weightMatrix_36_1),
    .io_weightMatrix_36_2(neuralNets_io_weightMatrix_36_2),
    .io_weightMatrix_36_3(neuralNets_io_weightMatrix_36_3),
    .io_weightMatrix_37_0(neuralNets_io_weightMatrix_37_0),
    .io_weightMatrix_37_1(neuralNets_io_weightMatrix_37_1),
    .io_weightMatrix_37_2(neuralNets_io_weightMatrix_37_2),
    .io_weightMatrix_37_3(neuralNets_io_weightMatrix_37_3),
    .io_weightMatrix_38_0(neuralNets_io_weightMatrix_38_0),
    .io_weightMatrix_38_1(neuralNets_io_weightMatrix_38_1),
    .io_weightMatrix_38_2(neuralNets_io_weightMatrix_38_2),
    .io_weightMatrix_38_3(neuralNets_io_weightMatrix_38_3),
    .io_weightMatrix_39_0(neuralNets_io_weightMatrix_39_0),
    .io_weightMatrix_39_1(neuralNets_io_weightMatrix_39_1),
    .io_weightMatrix_39_2(neuralNets_io_weightMatrix_39_2),
    .io_weightMatrix_39_3(neuralNets_io_weightMatrix_39_3),
    .io_weightMatrix_40_0(neuralNets_io_weightMatrix_40_0),
    .io_weightMatrix_40_1(neuralNets_io_weightMatrix_40_1),
    .io_weightMatrix_40_2(neuralNets_io_weightMatrix_40_2),
    .io_weightMatrix_40_3(neuralNets_io_weightMatrix_40_3),
    .io_weightMatrix_41_0(neuralNets_io_weightMatrix_41_0),
    .io_weightMatrix_41_1(neuralNets_io_weightMatrix_41_1),
    .io_weightMatrix_41_2(neuralNets_io_weightMatrix_41_2),
    .io_weightMatrix_41_3(neuralNets_io_weightMatrix_41_3),
    .io_weightMatrix_42_0(neuralNets_io_weightMatrix_42_0),
    .io_weightMatrix_42_1(neuralNets_io_weightMatrix_42_1),
    .io_weightMatrix_42_2(neuralNets_io_weightMatrix_42_2),
    .io_weightMatrix_42_3(neuralNets_io_weightMatrix_42_3),
    .io_weightMatrix_43_0(neuralNets_io_weightMatrix_43_0),
    .io_weightMatrix_43_1(neuralNets_io_weightMatrix_43_1),
    .io_weightMatrix_43_2(neuralNets_io_weightMatrix_43_2),
    .io_weightMatrix_43_3(neuralNets_io_weightMatrix_43_3),
    .io_weightMatrix_44_0(neuralNets_io_weightMatrix_44_0),
    .io_weightMatrix_44_1(neuralNets_io_weightMatrix_44_1),
    .io_weightMatrix_44_2(neuralNets_io_weightMatrix_44_2),
    .io_weightMatrix_44_3(neuralNets_io_weightMatrix_44_3),
    .io_weightMatrix_45_0(neuralNets_io_weightMatrix_45_0),
    .io_weightMatrix_45_1(neuralNets_io_weightMatrix_45_1),
    .io_weightMatrix_45_2(neuralNets_io_weightMatrix_45_2),
    .io_weightMatrix_45_3(neuralNets_io_weightMatrix_45_3),
    .io_weightMatrix_46_0(neuralNets_io_weightMatrix_46_0),
    .io_weightMatrix_46_1(neuralNets_io_weightMatrix_46_1),
    .io_weightMatrix_46_2(neuralNets_io_weightMatrix_46_2),
    .io_weightMatrix_46_3(neuralNets_io_weightMatrix_46_3),
    .io_weightMatrix_47_0(neuralNets_io_weightMatrix_47_0),
    .io_weightMatrix_47_1(neuralNets_io_weightMatrix_47_1),
    .io_weightMatrix_47_2(neuralNets_io_weightMatrix_47_2),
    .io_weightMatrix_47_3(neuralNets_io_weightMatrix_47_3),
    .io_weightMatrix_48_0(neuralNets_io_weightMatrix_48_0),
    .io_weightMatrix_48_1(neuralNets_io_weightMatrix_48_1),
    .io_weightMatrix_48_2(neuralNets_io_weightMatrix_48_2),
    .io_weightMatrix_48_3(neuralNets_io_weightMatrix_48_3),
    .io_weightMatrix_49_0(neuralNets_io_weightMatrix_49_0),
    .io_weightMatrix_49_1(neuralNets_io_weightMatrix_49_1),
    .io_weightMatrix_49_2(neuralNets_io_weightMatrix_49_2),
    .io_weightMatrix_49_3(neuralNets_io_weightMatrix_49_3),
    .io_weightMatrix_50_0(neuralNets_io_weightMatrix_50_0),
    .io_weightMatrix_50_1(neuralNets_io_weightMatrix_50_1),
    .io_weightMatrix_50_2(neuralNets_io_weightMatrix_50_2),
    .io_weightMatrix_50_3(neuralNets_io_weightMatrix_50_3),
    .io_weightMatrix_51_0(neuralNets_io_weightMatrix_51_0),
    .io_weightMatrix_51_1(neuralNets_io_weightMatrix_51_1),
    .io_weightMatrix_51_2(neuralNets_io_weightMatrix_51_2),
    .io_weightMatrix_51_3(neuralNets_io_weightMatrix_51_3),
    .io_weightMatrix_52_0(neuralNets_io_weightMatrix_52_0),
    .io_weightMatrix_52_1(neuralNets_io_weightMatrix_52_1),
    .io_weightMatrix_52_2(neuralNets_io_weightMatrix_52_2),
    .io_weightMatrix_52_3(neuralNets_io_weightMatrix_52_3),
    .io_weightMatrix_53_0(neuralNets_io_weightMatrix_53_0),
    .io_weightMatrix_53_1(neuralNets_io_weightMatrix_53_1),
    .io_weightMatrix_53_2(neuralNets_io_weightMatrix_53_2),
    .io_weightMatrix_53_3(neuralNets_io_weightMatrix_53_3),
    .io_weightMatrix_54_0(neuralNets_io_weightMatrix_54_0),
    .io_weightMatrix_54_1(neuralNets_io_weightMatrix_54_1),
    .io_weightMatrix_54_2(neuralNets_io_weightMatrix_54_2),
    .io_weightMatrix_54_3(neuralNets_io_weightMatrix_54_3),
    .io_weightMatrix_55_0(neuralNets_io_weightMatrix_55_0),
    .io_weightMatrix_55_1(neuralNets_io_weightMatrix_55_1),
    .io_weightMatrix_55_2(neuralNets_io_weightMatrix_55_2),
    .io_weightMatrix_55_3(neuralNets_io_weightMatrix_55_3),
    .io_weightMatrix_56_0(neuralNets_io_weightMatrix_56_0),
    .io_weightMatrix_56_1(neuralNets_io_weightMatrix_56_1),
    .io_weightMatrix_56_2(neuralNets_io_weightMatrix_56_2),
    .io_weightMatrix_56_3(neuralNets_io_weightMatrix_56_3),
    .io_weightMatrix_57_0(neuralNets_io_weightMatrix_57_0),
    .io_weightMatrix_57_1(neuralNets_io_weightMatrix_57_1),
    .io_weightMatrix_57_2(neuralNets_io_weightMatrix_57_2),
    .io_weightMatrix_57_3(neuralNets_io_weightMatrix_57_3),
    .io_weightMatrix_58_0(neuralNets_io_weightMatrix_58_0),
    .io_weightMatrix_58_1(neuralNets_io_weightMatrix_58_1),
    .io_weightMatrix_58_2(neuralNets_io_weightMatrix_58_2),
    .io_weightMatrix_58_3(neuralNets_io_weightMatrix_58_3),
    .io_weightMatrix_59_0(neuralNets_io_weightMatrix_59_0),
    .io_weightMatrix_59_1(neuralNets_io_weightMatrix_59_1),
    .io_weightMatrix_59_2(neuralNets_io_weightMatrix_59_2),
    .io_weightMatrix_59_3(neuralNets_io_weightMatrix_59_3),
    .io_weightMatrix_60_0(neuralNets_io_weightMatrix_60_0),
    .io_weightMatrix_60_1(neuralNets_io_weightMatrix_60_1),
    .io_weightMatrix_60_2(neuralNets_io_weightMatrix_60_2),
    .io_weightMatrix_60_3(neuralNets_io_weightMatrix_60_3),
    .io_weightMatrix_61_0(neuralNets_io_weightMatrix_61_0),
    .io_weightMatrix_61_1(neuralNets_io_weightMatrix_61_1),
    .io_weightMatrix_61_2(neuralNets_io_weightMatrix_61_2),
    .io_weightMatrix_61_3(neuralNets_io_weightMatrix_61_3),
    .io_weightMatrix_62_0(neuralNets_io_weightMatrix_62_0),
    .io_weightMatrix_62_1(neuralNets_io_weightMatrix_62_1),
    .io_weightMatrix_62_2(neuralNets_io_weightMatrix_62_2),
    .io_weightMatrix_62_3(neuralNets_io_weightMatrix_62_3),
    .io_weightMatrix_63_0(neuralNets_io_weightMatrix_63_0),
    .io_weightMatrix_63_1(neuralNets_io_weightMatrix_63_1),
    .io_weightMatrix_63_2(neuralNets_io_weightMatrix_63_2),
    .io_weightMatrix_63_3(neuralNets_io_weightMatrix_63_3),
    .io_weightMatrix_64_0(neuralNets_io_weightMatrix_64_0),
    .io_weightMatrix_64_1(neuralNets_io_weightMatrix_64_1),
    .io_weightMatrix_64_2(neuralNets_io_weightMatrix_64_2),
    .io_weightMatrix_64_3(neuralNets_io_weightMatrix_64_3),
    .io_weightMatrix_65_0(neuralNets_io_weightMatrix_65_0),
    .io_weightMatrix_65_1(neuralNets_io_weightMatrix_65_1),
    .io_weightMatrix_65_2(neuralNets_io_weightMatrix_65_2),
    .io_weightMatrix_65_3(neuralNets_io_weightMatrix_65_3),
    .io_weightMatrix_66_0(neuralNets_io_weightMatrix_66_0),
    .io_weightMatrix_66_1(neuralNets_io_weightMatrix_66_1),
    .io_weightMatrix_66_2(neuralNets_io_weightMatrix_66_2),
    .io_weightMatrix_66_3(neuralNets_io_weightMatrix_66_3),
    .io_weightMatrix_67_0(neuralNets_io_weightMatrix_67_0),
    .io_weightMatrix_67_1(neuralNets_io_weightMatrix_67_1),
    .io_weightMatrix_67_2(neuralNets_io_weightMatrix_67_2),
    .io_weightMatrix_67_3(neuralNets_io_weightMatrix_67_3),
    .io_weightMatrix_68_0(neuralNets_io_weightMatrix_68_0),
    .io_weightMatrix_68_1(neuralNets_io_weightMatrix_68_1),
    .io_weightMatrix_68_2(neuralNets_io_weightMatrix_68_2),
    .io_weightMatrix_68_3(neuralNets_io_weightMatrix_68_3),
    .io_weightMatrix_69_0(neuralNets_io_weightMatrix_69_0),
    .io_weightMatrix_69_1(neuralNets_io_weightMatrix_69_1),
    .io_weightMatrix_69_2(neuralNets_io_weightMatrix_69_2),
    .io_weightMatrix_69_3(neuralNets_io_weightMatrix_69_3),
    .io_weightMatrix_70_0(neuralNets_io_weightMatrix_70_0),
    .io_weightMatrix_70_1(neuralNets_io_weightMatrix_70_1),
    .io_weightMatrix_70_2(neuralNets_io_weightMatrix_70_2),
    .io_weightMatrix_70_3(neuralNets_io_weightMatrix_70_3),
    .io_weightMatrix_71_0(neuralNets_io_weightMatrix_71_0),
    .io_weightMatrix_71_1(neuralNets_io_weightMatrix_71_1),
    .io_weightMatrix_71_2(neuralNets_io_weightMatrix_71_2),
    .io_weightMatrix_71_3(neuralNets_io_weightMatrix_71_3),
    .io_weightMatrix_72_0(neuralNets_io_weightMatrix_72_0),
    .io_weightMatrix_72_1(neuralNets_io_weightMatrix_72_1),
    .io_weightMatrix_72_2(neuralNets_io_weightMatrix_72_2),
    .io_weightMatrix_72_3(neuralNets_io_weightMatrix_72_3),
    .io_weightMatrix_73_0(neuralNets_io_weightMatrix_73_0),
    .io_weightMatrix_73_1(neuralNets_io_weightMatrix_73_1),
    .io_weightMatrix_73_2(neuralNets_io_weightMatrix_73_2),
    .io_weightMatrix_73_3(neuralNets_io_weightMatrix_73_3),
    .io_weightMatrix_74_0(neuralNets_io_weightMatrix_74_0),
    .io_weightMatrix_74_1(neuralNets_io_weightMatrix_74_1),
    .io_weightMatrix_74_2(neuralNets_io_weightMatrix_74_2),
    .io_weightMatrix_74_3(neuralNets_io_weightMatrix_74_3),
    .io_weightMatrix_75_0(neuralNets_io_weightMatrix_75_0),
    .io_weightMatrix_75_1(neuralNets_io_weightMatrix_75_1),
    .io_weightMatrix_75_2(neuralNets_io_weightMatrix_75_2),
    .io_weightMatrix_75_3(neuralNets_io_weightMatrix_75_3),
    .io_weightMatrix_76_0(neuralNets_io_weightMatrix_76_0),
    .io_weightMatrix_76_1(neuralNets_io_weightMatrix_76_1),
    .io_weightMatrix_76_2(neuralNets_io_weightMatrix_76_2),
    .io_weightMatrix_76_3(neuralNets_io_weightMatrix_76_3),
    .io_weightMatrix_77_0(neuralNets_io_weightMatrix_77_0),
    .io_weightMatrix_77_1(neuralNets_io_weightMatrix_77_1),
    .io_weightMatrix_77_2(neuralNets_io_weightMatrix_77_2),
    .io_weightMatrix_77_3(neuralNets_io_weightMatrix_77_3),
    .io_weightMatrix_78_0(neuralNets_io_weightMatrix_78_0),
    .io_weightMatrix_78_1(neuralNets_io_weightMatrix_78_1),
    .io_weightMatrix_78_2(neuralNets_io_weightMatrix_78_2),
    .io_weightMatrix_78_3(neuralNets_io_weightMatrix_78_3),
    .io_weightMatrix_79_0(neuralNets_io_weightMatrix_79_0),
    .io_weightMatrix_79_1(neuralNets_io_weightMatrix_79_1),
    .io_weightMatrix_79_2(neuralNets_io_weightMatrix_79_2),
    .io_weightMatrix_79_3(neuralNets_io_weightMatrix_79_3),
    .io_weightMatrix_80_0(neuralNets_io_weightMatrix_80_0),
    .io_weightMatrix_80_1(neuralNets_io_weightMatrix_80_1),
    .io_weightMatrix_80_2(neuralNets_io_weightMatrix_80_2),
    .io_weightMatrix_80_3(neuralNets_io_weightMatrix_80_3),
    .io_weightMatrix_81_0(neuralNets_io_weightMatrix_81_0),
    .io_weightMatrix_81_1(neuralNets_io_weightMatrix_81_1),
    .io_weightMatrix_81_2(neuralNets_io_weightMatrix_81_2),
    .io_weightMatrix_81_3(neuralNets_io_weightMatrix_81_3),
    .io_weightMatrix_82_0(neuralNets_io_weightMatrix_82_0),
    .io_weightMatrix_82_1(neuralNets_io_weightMatrix_82_1),
    .io_weightMatrix_82_2(neuralNets_io_weightMatrix_82_2),
    .io_weightMatrix_82_3(neuralNets_io_weightMatrix_82_3),
    .io_weightMatrix_83_0(neuralNets_io_weightMatrix_83_0),
    .io_weightMatrix_83_1(neuralNets_io_weightMatrix_83_1),
    .io_weightMatrix_83_2(neuralNets_io_weightMatrix_83_2),
    .io_weightMatrix_83_3(neuralNets_io_weightMatrix_83_3),
    .io_weightMatrix_84_0(neuralNets_io_weightMatrix_84_0),
    .io_weightMatrix_84_1(neuralNets_io_weightMatrix_84_1),
    .io_weightMatrix_84_2(neuralNets_io_weightMatrix_84_2),
    .io_weightMatrix_84_3(neuralNets_io_weightMatrix_84_3),
    .io_weightMatrix_85_0(neuralNets_io_weightMatrix_85_0),
    .io_weightMatrix_85_1(neuralNets_io_weightMatrix_85_1),
    .io_weightMatrix_85_2(neuralNets_io_weightMatrix_85_2),
    .io_weightMatrix_85_3(neuralNets_io_weightMatrix_85_3),
    .io_weightMatrix_86_0(neuralNets_io_weightMatrix_86_0),
    .io_weightMatrix_86_1(neuralNets_io_weightMatrix_86_1),
    .io_weightMatrix_86_2(neuralNets_io_weightMatrix_86_2),
    .io_weightMatrix_86_3(neuralNets_io_weightMatrix_86_3),
    .io_weightMatrix_87_0(neuralNets_io_weightMatrix_87_0),
    .io_weightMatrix_87_1(neuralNets_io_weightMatrix_87_1),
    .io_weightMatrix_87_2(neuralNets_io_weightMatrix_87_2),
    .io_weightMatrix_87_3(neuralNets_io_weightMatrix_87_3),
    .io_weightMatrix_88_0(neuralNets_io_weightMatrix_88_0),
    .io_weightMatrix_88_1(neuralNets_io_weightMatrix_88_1),
    .io_weightMatrix_88_2(neuralNets_io_weightMatrix_88_2),
    .io_weightMatrix_88_3(neuralNets_io_weightMatrix_88_3),
    .io_weightMatrix_89_0(neuralNets_io_weightMatrix_89_0),
    .io_weightMatrix_89_1(neuralNets_io_weightMatrix_89_1),
    .io_weightMatrix_89_2(neuralNets_io_weightMatrix_89_2),
    .io_weightMatrix_89_3(neuralNets_io_weightMatrix_89_3),
    .io_weightMatrix_90_0(neuralNets_io_weightMatrix_90_0),
    .io_weightMatrix_90_1(neuralNets_io_weightMatrix_90_1),
    .io_weightMatrix_90_2(neuralNets_io_weightMatrix_90_2),
    .io_weightMatrix_90_3(neuralNets_io_weightMatrix_90_3),
    .io_weightMatrix_91_0(neuralNets_io_weightMatrix_91_0),
    .io_weightMatrix_91_1(neuralNets_io_weightMatrix_91_1),
    .io_weightMatrix_91_2(neuralNets_io_weightMatrix_91_2),
    .io_weightMatrix_91_3(neuralNets_io_weightMatrix_91_3),
    .io_weightMatrix_92_0(neuralNets_io_weightMatrix_92_0),
    .io_weightMatrix_92_1(neuralNets_io_weightMatrix_92_1),
    .io_weightMatrix_92_2(neuralNets_io_weightMatrix_92_2),
    .io_weightMatrix_92_3(neuralNets_io_weightMatrix_92_3),
    .io_weightMatrix_93_0(neuralNets_io_weightMatrix_93_0),
    .io_weightMatrix_93_1(neuralNets_io_weightMatrix_93_1),
    .io_weightMatrix_93_2(neuralNets_io_weightMatrix_93_2),
    .io_weightMatrix_93_3(neuralNets_io_weightMatrix_93_3),
    .io_weightMatrix_94_0(neuralNets_io_weightMatrix_94_0),
    .io_weightMatrix_94_1(neuralNets_io_weightMatrix_94_1),
    .io_weightMatrix_94_2(neuralNets_io_weightMatrix_94_2),
    .io_weightMatrix_94_3(neuralNets_io_weightMatrix_94_3),
    .io_weightMatrix_95_0(neuralNets_io_weightMatrix_95_0),
    .io_weightMatrix_95_1(neuralNets_io_weightMatrix_95_1),
    .io_weightMatrix_95_2(neuralNets_io_weightMatrix_95_2),
    .io_weightMatrix_95_3(neuralNets_io_weightMatrix_95_3),
    .io_weightMatrix_96_0(neuralNets_io_weightMatrix_96_0),
    .io_weightMatrix_96_1(neuralNets_io_weightMatrix_96_1),
    .io_weightMatrix_96_2(neuralNets_io_weightMatrix_96_2),
    .io_weightMatrix_96_3(neuralNets_io_weightMatrix_96_3),
    .io_weightMatrix_97_0(neuralNets_io_weightMatrix_97_0),
    .io_weightMatrix_97_1(neuralNets_io_weightMatrix_97_1),
    .io_weightMatrix_97_2(neuralNets_io_weightMatrix_97_2),
    .io_weightMatrix_97_3(neuralNets_io_weightMatrix_97_3),
    .io_weightMatrix_98_0(neuralNets_io_weightMatrix_98_0),
    .io_weightMatrix_98_1(neuralNets_io_weightMatrix_98_1),
    .io_weightMatrix_98_2(neuralNets_io_weightMatrix_98_2),
    .io_weightMatrix_98_3(neuralNets_io_weightMatrix_98_3),
    .io_weightMatrix_99_0(neuralNets_io_weightMatrix_99_0),
    .io_weightMatrix_99_1(neuralNets_io_weightMatrix_99_1),
    .io_weightMatrix_99_2(neuralNets_io_weightMatrix_99_2),
    .io_weightMatrix_99_3(neuralNets_io_weightMatrix_99_3),
    .io_weightVec_0(neuralNets_io_weightVec_0),
    .io_weightVec_1(neuralNets_io_weightVec_1),
    .io_weightVec_2(neuralNets_io_weightVec_2),
    .io_weightVec_3(neuralNets_io_weightVec_3),
    .io_weightVec_4(neuralNets_io_weightVec_4),
    .io_weightVec_5(neuralNets_io_weightVec_5),
    .io_weightVec_6(neuralNets_io_weightVec_6),
    .io_weightVec_7(neuralNets_io_weightVec_7),
    .io_weightVec_8(neuralNets_io_weightVec_8),
    .io_weightVec_9(neuralNets_io_weightVec_9),
    .io_weightVec_10(neuralNets_io_weightVec_10),
    .io_weightVec_11(neuralNets_io_weightVec_11),
    .io_weightVec_12(neuralNets_io_weightVec_12),
    .io_weightVec_13(neuralNets_io_weightVec_13),
    .io_weightVec_14(neuralNets_io_weightVec_14),
    .io_weightVec_15(neuralNets_io_weightVec_15),
    .io_weightVec_16(neuralNets_io_weightVec_16),
    .io_weightVec_17(neuralNets_io_weightVec_17),
    .io_weightVec_18(neuralNets_io_weightVec_18),
    .io_weightVec_19(neuralNets_io_weightVec_19),
    .io_weightVec_20(neuralNets_io_weightVec_20),
    .io_weightVec_21(neuralNets_io_weightVec_21),
    .io_weightVec_22(neuralNets_io_weightVec_22),
    .io_weightVec_23(neuralNets_io_weightVec_23),
    .io_weightVec_24(neuralNets_io_weightVec_24),
    .io_weightVec_25(neuralNets_io_weightVec_25),
    .io_weightVec_26(neuralNets_io_weightVec_26),
    .io_weightVec_27(neuralNets_io_weightVec_27),
    .io_weightVec_28(neuralNets_io_weightVec_28),
    .io_weightVec_29(neuralNets_io_weightVec_29),
    .io_weightVec_30(neuralNets_io_weightVec_30),
    .io_weightVec_31(neuralNets_io_weightVec_31),
    .io_weightVec_32(neuralNets_io_weightVec_32),
    .io_weightVec_33(neuralNets_io_weightVec_33),
    .io_weightVec_34(neuralNets_io_weightVec_34),
    .io_weightVec_35(neuralNets_io_weightVec_35),
    .io_weightVec_36(neuralNets_io_weightVec_36),
    .io_weightVec_37(neuralNets_io_weightVec_37),
    .io_weightVec_38(neuralNets_io_weightVec_38),
    .io_weightVec_39(neuralNets_io_weightVec_39),
    .io_weightVec_40(neuralNets_io_weightVec_40),
    .io_weightVec_41(neuralNets_io_weightVec_41),
    .io_weightVec_42(neuralNets_io_weightVec_42),
    .io_weightVec_43(neuralNets_io_weightVec_43),
    .io_weightVec_44(neuralNets_io_weightVec_44),
    .io_weightVec_45(neuralNets_io_weightVec_45),
    .io_weightVec_46(neuralNets_io_weightVec_46),
    .io_weightVec_47(neuralNets_io_weightVec_47),
    .io_weightVec_48(neuralNets_io_weightVec_48),
    .io_weightVec_49(neuralNets_io_weightVec_49),
    .io_weightVec_50(neuralNets_io_weightVec_50),
    .io_weightVec_51(neuralNets_io_weightVec_51),
    .io_weightVec_52(neuralNets_io_weightVec_52),
    .io_weightVec_53(neuralNets_io_weightVec_53),
    .io_weightVec_54(neuralNets_io_weightVec_54),
    .io_weightVec_55(neuralNets_io_weightVec_55),
    .io_weightVec_56(neuralNets_io_weightVec_56),
    .io_weightVec_57(neuralNets_io_weightVec_57),
    .io_weightVec_58(neuralNets_io_weightVec_58),
    .io_weightVec_59(neuralNets_io_weightVec_59),
    .io_weightVec_60(neuralNets_io_weightVec_60),
    .io_weightVec_61(neuralNets_io_weightVec_61),
    .io_weightVec_62(neuralNets_io_weightVec_62),
    .io_weightVec_63(neuralNets_io_weightVec_63),
    .io_weightVec_64(neuralNets_io_weightVec_64),
    .io_weightVec_65(neuralNets_io_weightVec_65),
    .io_weightVec_66(neuralNets_io_weightVec_66),
    .io_weightVec_67(neuralNets_io_weightVec_67),
    .io_weightVec_68(neuralNets_io_weightVec_68),
    .io_weightVec_69(neuralNets_io_weightVec_69),
    .io_weightVec_70(neuralNets_io_weightVec_70),
    .io_weightVec_71(neuralNets_io_weightVec_71),
    .io_weightVec_72(neuralNets_io_weightVec_72),
    .io_weightVec_73(neuralNets_io_weightVec_73),
    .io_weightVec_74(neuralNets_io_weightVec_74),
    .io_weightVec_75(neuralNets_io_weightVec_75),
    .io_weightVec_76(neuralNets_io_weightVec_76),
    .io_weightVec_77(neuralNets_io_weightVec_77),
    .io_weightVec_78(neuralNets_io_weightVec_78),
    .io_weightVec_79(neuralNets_io_weightVec_79),
    .io_weightVec_80(neuralNets_io_weightVec_80),
    .io_weightVec_81(neuralNets_io_weightVec_81),
    .io_weightVec_82(neuralNets_io_weightVec_82),
    .io_weightVec_83(neuralNets_io_weightVec_83),
    .io_weightVec_84(neuralNets_io_weightVec_84),
    .io_weightVec_85(neuralNets_io_weightVec_85),
    .io_weightVec_86(neuralNets_io_weightVec_86),
    .io_weightVec_87(neuralNets_io_weightVec_87),
    .io_weightVec_88(neuralNets_io_weightVec_88),
    .io_weightVec_89(neuralNets_io_weightVec_89),
    .io_weightVec_90(neuralNets_io_weightVec_90),
    .io_weightVec_91(neuralNets_io_weightVec_91),
    .io_weightVec_92(neuralNets_io_weightVec_92),
    .io_weightVec_93(neuralNets_io_weightVec_93),
    .io_weightVec_94(neuralNets_io_weightVec_94),
    .io_weightVec_95(neuralNets_io_weightVec_95),
    .io_weightVec_96(neuralNets_io_weightVec_96),
    .io_weightVec_97(neuralNets_io_weightVec_97),
    .io_weightVec_98(neuralNets_io_weightVec_98),
    .io_weightVec_99(neuralNets_io_weightVec_99),
    .io_biasVec_0(neuralNets_io_biasVec_0),
    .io_biasVec_1(neuralNets_io_biasVec_1),
    .io_biasVec_2(neuralNets_io_biasVec_2),
    .io_biasVec_3(neuralNets_io_biasVec_3),
    .io_biasVec_4(neuralNets_io_biasVec_4),
    .io_biasVec_5(neuralNets_io_biasVec_5),
    .io_biasVec_6(neuralNets_io_biasVec_6),
    .io_biasVec_7(neuralNets_io_biasVec_7),
    .io_biasVec_8(neuralNets_io_biasVec_8),
    .io_biasVec_9(neuralNets_io_biasVec_9),
    .io_biasVec_10(neuralNets_io_biasVec_10),
    .io_biasVec_11(neuralNets_io_biasVec_11),
    .io_biasVec_12(neuralNets_io_biasVec_12),
    .io_biasVec_13(neuralNets_io_biasVec_13),
    .io_biasVec_14(neuralNets_io_biasVec_14),
    .io_biasVec_15(neuralNets_io_biasVec_15),
    .io_biasVec_16(neuralNets_io_biasVec_16),
    .io_biasVec_17(neuralNets_io_biasVec_17),
    .io_biasVec_18(neuralNets_io_biasVec_18),
    .io_biasVec_19(neuralNets_io_biasVec_19),
    .io_biasVec_20(neuralNets_io_biasVec_20),
    .io_biasVec_21(neuralNets_io_biasVec_21),
    .io_biasVec_22(neuralNets_io_biasVec_22),
    .io_biasVec_23(neuralNets_io_biasVec_23),
    .io_biasVec_24(neuralNets_io_biasVec_24),
    .io_biasVec_25(neuralNets_io_biasVec_25),
    .io_biasVec_26(neuralNets_io_biasVec_26),
    .io_biasVec_27(neuralNets_io_biasVec_27),
    .io_biasVec_28(neuralNets_io_biasVec_28),
    .io_biasVec_29(neuralNets_io_biasVec_29),
    .io_biasVec_30(neuralNets_io_biasVec_30),
    .io_biasVec_31(neuralNets_io_biasVec_31),
    .io_biasVec_32(neuralNets_io_biasVec_32),
    .io_biasVec_33(neuralNets_io_biasVec_33),
    .io_biasVec_34(neuralNets_io_biasVec_34),
    .io_biasVec_35(neuralNets_io_biasVec_35),
    .io_biasVec_36(neuralNets_io_biasVec_36),
    .io_biasVec_37(neuralNets_io_biasVec_37),
    .io_biasVec_38(neuralNets_io_biasVec_38),
    .io_biasVec_39(neuralNets_io_biasVec_39),
    .io_biasVec_40(neuralNets_io_biasVec_40),
    .io_biasVec_41(neuralNets_io_biasVec_41),
    .io_biasVec_42(neuralNets_io_biasVec_42),
    .io_biasVec_43(neuralNets_io_biasVec_43),
    .io_biasVec_44(neuralNets_io_biasVec_44),
    .io_biasVec_45(neuralNets_io_biasVec_45),
    .io_biasVec_46(neuralNets_io_biasVec_46),
    .io_biasVec_47(neuralNets_io_biasVec_47),
    .io_biasVec_48(neuralNets_io_biasVec_48),
    .io_biasVec_49(neuralNets_io_biasVec_49),
    .io_biasVec_50(neuralNets_io_biasVec_50),
    .io_biasVec_51(neuralNets_io_biasVec_51),
    .io_biasVec_52(neuralNets_io_biasVec_52),
    .io_biasVec_53(neuralNets_io_biasVec_53),
    .io_biasVec_54(neuralNets_io_biasVec_54),
    .io_biasVec_55(neuralNets_io_biasVec_55),
    .io_biasVec_56(neuralNets_io_biasVec_56),
    .io_biasVec_57(neuralNets_io_biasVec_57),
    .io_biasVec_58(neuralNets_io_biasVec_58),
    .io_biasVec_59(neuralNets_io_biasVec_59),
    .io_biasVec_60(neuralNets_io_biasVec_60),
    .io_biasVec_61(neuralNets_io_biasVec_61),
    .io_biasVec_62(neuralNets_io_biasVec_62),
    .io_biasVec_63(neuralNets_io_biasVec_63),
    .io_biasVec_64(neuralNets_io_biasVec_64),
    .io_biasVec_65(neuralNets_io_biasVec_65),
    .io_biasVec_66(neuralNets_io_biasVec_66),
    .io_biasVec_67(neuralNets_io_biasVec_67),
    .io_biasVec_68(neuralNets_io_biasVec_68),
    .io_biasVec_69(neuralNets_io_biasVec_69),
    .io_biasVec_70(neuralNets_io_biasVec_70),
    .io_biasVec_71(neuralNets_io_biasVec_71),
    .io_biasVec_72(neuralNets_io_biasVec_72),
    .io_biasVec_73(neuralNets_io_biasVec_73),
    .io_biasVec_74(neuralNets_io_biasVec_74),
    .io_biasVec_75(neuralNets_io_biasVec_75),
    .io_biasVec_76(neuralNets_io_biasVec_76),
    .io_biasVec_77(neuralNets_io_biasVec_77),
    .io_biasVec_78(neuralNets_io_biasVec_78),
    .io_biasVec_79(neuralNets_io_biasVec_79),
    .io_biasVec_80(neuralNets_io_biasVec_80),
    .io_biasVec_81(neuralNets_io_biasVec_81),
    .io_biasVec_82(neuralNets_io_biasVec_82),
    .io_biasVec_83(neuralNets_io_biasVec_83),
    .io_biasVec_84(neuralNets_io_biasVec_84),
    .io_biasVec_85(neuralNets_io_biasVec_85),
    .io_biasVec_86(neuralNets_io_biasVec_86),
    .io_biasVec_87(neuralNets_io_biasVec_87),
    .io_biasVec_88(neuralNets_io_biasVec_88),
    .io_biasVec_89(neuralNets_io_biasVec_89),
    .io_biasVec_90(neuralNets_io_biasVec_90),
    .io_biasVec_91(neuralNets_io_biasVec_91),
    .io_biasVec_92(neuralNets_io_biasVec_92),
    .io_biasVec_93(neuralNets_io_biasVec_93),
    .io_biasVec_94(neuralNets_io_biasVec_94),
    .io_biasVec_95(neuralNets_io_biasVec_95),
    .io_biasVec_96(neuralNets_io_biasVec_96),
    .io_biasVec_97(neuralNets_io_biasVec_97),
    .io_biasVec_98(neuralNets_io_biasVec_98),
    .io_biasVec_99(neuralNets_io_biasVec_99),
    .io_biasScalar(neuralNets_io_biasScalar),
    .io_rawVotes(neuralNets_io_rawVotes)
  );
  assign _T_1 = $unsigned(io_streamIn_bits); // @[Wellness.scala 271:80]
  assign _T_2 = $signed(_T_1); // @[Wellness.scala 271:80]
  assign _T_4 = $unsigned(io_in_bits); // @[Wellness.scala 271:125]
  assign _T_5 = $signed(_T_4); // @[Wellness.scala 271:125]
  assign _T_10 = $unsigned(filter1_io_out_bits); // @[Wellness.scala 283:57]
  assign _T_22 = $unsigned(lineLength1_io_out_bits); // @[Wellness.scala 314:65]
  assign _T_25 = $unsigned(bandpowerAlpha_io_out_bits); // @[Wellness.scala 327:58]
  assign _T_28 = $unsigned(bandpowerBeta_io_out_bits); // @[Wellness.scala 328:57]
  assign _T_31 = $unsigned(bandpowerGamma_io_out_bits); // @[Wellness.scala 329:58]
  assign _T_34 = $unsigned(lineLength1Reg1); // @[Wellness.scala 330:47]
  assign _T_36 = lineLength1Valid1 & bandpowerAlpha_io_out_valid; // @[Wellness.scala 332:48]
  assign _T_37 = _T_36 & bandpowerBeta_io_out_valid; // @[Wellness.scala 332:79]
  assign io_out_valid = neuralNets_io_out_valid; // @[Wellness.scala 342:16]
  assign io_out_bits = neuralNets_io_out_bits; // @[Wellness.scala 344:15]
  assign io_rawVotes = neuralNets_io_rawVotes; // @[Wellness.scala 345:15]
  assign filter1_clock = clock;
  assign filter1_reset = reset;
  assign filter1_io_in_valid = io_inConf_bits_confInputMuxSel ? io_streamIn_valid : io_in_valid; // @[Wellness.scala 276:23]
  assign filter1_io_in_bits = io_inConf_bits_confInputMuxSel ? $signed(_T_2) : $signed(_T_5); // @[Wellness.scala 278:22]
  assign lineLength1_clock = clock;
  assign lineLength1_reset = reset;
  assign lineLength1_io_in_valid = filter1_io_out_valid; // @[Wellness.scala 281:27]
  assign lineLength1_io_in_bits = $signed(_T_10); // @[Wellness.scala 283:26]
  assign filterAlpha_clock = clock;
  assign filterAlpha_reset = reset;
  assign filterAlpha_io_in_valid = filter1_io_out_valid; // @[Wellness.scala 286:27]
  assign filterAlpha_io_in_bits = $signed(_T_10); // @[Wellness.scala 288:26]
  assign filterBeta_clock = clock;
  assign filterBeta_reset = reset;
  assign filterBeta_io_in_valid = filter1_io_out_valid; // @[Wellness.scala 290:26]
  assign filterBeta_io_in_bits = $signed(_T_10); // @[Wellness.scala 292:25]
  assign filterGamma_clock = clock;
  assign filterGamma_reset = reset;
  assign filterGamma_io_in_valid = filter1_io_out_valid; // @[Wellness.scala 294:27]
  assign filterGamma_io_in_bits = $signed(_T_10); // @[Wellness.scala 296:26]
  assign bandpowerAlpha_clock = clock;
  assign bandpowerAlpha_reset = reset;
  assign bandpowerAlpha_io_in_valid = filterAlpha_io_out_valid; // @[Wellness.scala 300:30]
  assign bandpowerAlpha_io_in_bits = filterAlpha_io_out_bits; // @[Wellness.scala 302:29]
  assign bandpowerBeta_clock = clock;
  assign bandpowerBeta_reset = reset;
  assign bandpowerBeta_io_in_valid = filterBeta_io_out_valid; // @[Wellness.scala 304:29]
  assign bandpowerBeta_io_in_bits = filterBeta_io_out_bits; // @[Wellness.scala 306:28]
  assign bandpowerGamma_clock = clock;
  assign bandpowerGamma_reset = reset;
  assign bandpowerGamma_io_in_valid = filterGamma_io_out_valid; // @[Wellness.scala 308:30]
  assign bandpowerGamma_io_in_bits = filterGamma_io_out_bits; // @[Wellness.scala 310:29]
  assign neuralNets_clock = clock;
  assign neuralNets_io_in_valid = _T_37 & bandpowerGamma_io_out_valid; // @[Wellness.scala 332:26]
  assign neuralNets_io_in_bits_0 = $signed(_T_25); // @[Wellness.scala 333:25]
  assign neuralNets_io_in_bits_1 = $signed(_T_28); // @[Wellness.scala 333:25]
  assign neuralNets_io_in_bits_2 = $signed(_T_31); // @[Wellness.scala 333:25]
  assign neuralNets_io_in_bits_3 = $signed(_T_34); // @[Wellness.scala 333:25]
  assign neuralNets_io_weightMatrix_0_0 = io_inConf_bits_confneuralNetsweightMatrix_0_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_0_1 = io_inConf_bits_confneuralNetsweightMatrix_0_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_0_2 = io_inConf_bits_confneuralNetsweightMatrix_0_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_0_3 = io_inConf_bits_confneuralNetsweightMatrix_0_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_1_0 = io_inConf_bits_confneuralNetsweightMatrix_1_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_1_1 = io_inConf_bits_confneuralNetsweightMatrix_1_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_1_2 = io_inConf_bits_confneuralNetsweightMatrix_1_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_1_3 = io_inConf_bits_confneuralNetsweightMatrix_1_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_2_0 = io_inConf_bits_confneuralNetsweightMatrix_2_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_2_1 = io_inConf_bits_confneuralNetsweightMatrix_2_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_2_2 = io_inConf_bits_confneuralNetsweightMatrix_2_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_2_3 = io_inConf_bits_confneuralNetsweightMatrix_2_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_3_0 = io_inConf_bits_confneuralNetsweightMatrix_3_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_3_1 = io_inConf_bits_confneuralNetsweightMatrix_3_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_3_2 = io_inConf_bits_confneuralNetsweightMatrix_3_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_3_3 = io_inConf_bits_confneuralNetsweightMatrix_3_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_4_0 = io_inConf_bits_confneuralNetsweightMatrix_4_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_4_1 = io_inConf_bits_confneuralNetsweightMatrix_4_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_4_2 = io_inConf_bits_confneuralNetsweightMatrix_4_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_4_3 = io_inConf_bits_confneuralNetsweightMatrix_4_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_5_0 = io_inConf_bits_confneuralNetsweightMatrix_5_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_5_1 = io_inConf_bits_confneuralNetsweightMatrix_5_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_5_2 = io_inConf_bits_confneuralNetsweightMatrix_5_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_5_3 = io_inConf_bits_confneuralNetsweightMatrix_5_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_6_0 = io_inConf_bits_confneuralNetsweightMatrix_6_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_6_1 = io_inConf_bits_confneuralNetsweightMatrix_6_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_6_2 = io_inConf_bits_confneuralNetsweightMatrix_6_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_6_3 = io_inConf_bits_confneuralNetsweightMatrix_6_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_7_0 = io_inConf_bits_confneuralNetsweightMatrix_7_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_7_1 = io_inConf_bits_confneuralNetsweightMatrix_7_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_7_2 = io_inConf_bits_confneuralNetsweightMatrix_7_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_7_3 = io_inConf_bits_confneuralNetsweightMatrix_7_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_8_0 = io_inConf_bits_confneuralNetsweightMatrix_8_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_8_1 = io_inConf_bits_confneuralNetsweightMatrix_8_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_8_2 = io_inConf_bits_confneuralNetsweightMatrix_8_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_8_3 = io_inConf_bits_confneuralNetsweightMatrix_8_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_9_0 = io_inConf_bits_confneuralNetsweightMatrix_9_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_9_1 = io_inConf_bits_confneuralNetsweightMatrix_9_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_9_2 = io_inConf_bits_confneuralNetsweightMatrix_9_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_9_3 = io_inConf_bits_confneuralNetsweightMatrix_9_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_10_0 = io_inConf_bits_confneuralNetsweightMatrix_10_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_10_1 = io_inConf_bits_confneuralNetsweightMatrix_10_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_10_2 = io_inConf_bits_confneuralNetsweightMatrix_10_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_10_3 = io_inConf_bits_confneuralNetsweightMatrix_10_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_11_0 = io_inConf_bits_confneuralNetsweightMatrix_11_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_11_1 = io_inConf_bits_confneuralNetsweightMatrix_11_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_11_2 = io_inConf_bits_confneuralNetsweightMatrix_11_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_11_3 = io_inConf_bits_confneuralNetsweightMatrix_11_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_12_0 = io_inConf_bits_confneuralNetsweightMatrix_12_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_12_1 = io_inConf_bits_confneuralNetsweightMatrix_12_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_12_2 = io_inConf_bits_confneuralNetsweightMatrix_12_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_12_3 = io_inConf_bits_confneuralNetsweightMatrix_12_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_13_0 = io_inConf_bits_confneuralNetsweightMatrix_13_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_13_1 = io_inConf_bits_confneuralNetsweightMatrix_13_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_13_2 = io_inConf_bits_confneuralNetsweightMatrix_13_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_13_3 = io_inConf_bits_confneuralNetsweightMatrix_13_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_14_0 = io_inConf_bits_confneuralNetsweightMatrix_14_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_14_1 = io_inConf_bits_confneuralNetsweightMatrix_14_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_14_2 = io_inConf_bits_confneuralNetsweightMatrix_14_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_14_3 = io_inConf_bits_confneuralNetsweightMatrix_14_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_15_0 = io_inConf_bits_confneuralNetsweightMatrix_15_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_15_1 = io_inConf_bits_confneuralNetsweightMatrix_15_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_15_2 = io_inConf_bits_confneuralNetsweightMatrix_15_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_15_3 = io_inConf_bits_confneuralNetsweightMatrix_15_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_16_0 = io_inConf_bits_confneuralNetsweightMatrix_16_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_16_1 = io_inConf_bits_confneuralNetsweightMatrix_16_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_16_2 = io_inConf_bits_confneuralNetsweightMatrix_16_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_16_3 = io_inConf_bits_confneuralNetsweightMatrix_16_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_17_0 = io_inConf_bits_confneuralNetsweightMatrix_17_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_17_1 = io_inConf_bits_confneuralNetsweightMatrix_17_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_17_2 = io_inConf_bits_confneuralNetsweightMatrix_17_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_17_3 = io_inConf_bits_confneuralNetsweightMatrix_17_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_18_0 = io_inConf_bits_confneuralNetsweightMatrix_18_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_18_1 = io_inConf_bits_confneuralNetsweightMatrix_18_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_18_2 = io_inConf_bits_confneuralNetsweightMatrix_18_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_18_3 = io_inConf_bits_confneuralNetsweightMatrix_18_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_19_0 = io_inConf_bits_confneuralNetsweightMatrix_19_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_19_1 = io_inConf_bits_confneuralNetsweightMatrix_19_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_19_2 = io_inConf_bits_confneuralNetsweightMatrix_19_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_19_3 = io_inConf_bits_confneuralNetsweightMatrix_19_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_20_0 = io_inConf_bits_confneuralNetsweightMatrix_20_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_20_1 = io_inConf_bits_confneuralNetsweightMatrix_20_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_20_2 = io_inConf_bits_confneuralNetsweightMatrix_20_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_20_3 = io_inConf_bits_confneuralNetsweightMatrix_20_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_21_0 = io_inConf_bits_confneuralNetsweightMatrix_21_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_21_1 = io_inConf_bits_confneuralNetsweightMatrix_21_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_21_2 = io_inConf_bits_confneuralNetsweightMatrix_21_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_21_3 = io_inConf_bits_confneuralNetsweightMatrix_21_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_22_0 = io_inConf_bits_confneuralNetsweightMatrix_22_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_22_1 = io_inConf_bits_confneuralNetsweightMatrix_22_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_22_2 = io_inConf_bits_confneuralNetsweightMatrix_22_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_22_3 = io_inConf_bits_confneuralNetsweightMatrix_22_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_23_0 = io_inConf_bits_confneuralNetsweightMatrix_23_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_23_1 = io_inConf_bits_confneuralNetsweightMatrix_23_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_23_2 = io_inConf_bits_confneuralNetsweightMatrix_23_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_23_3 = io_inConf_bits_confneuralNetsweightMatrix_23_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_24_0 = io_inConf_bits_confneuralNetsweightMatrix_24_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_24_1 = io_inConf_bits_confneuralNetsweightMatrix_24_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_24_2 = io_inConf_bits_confneuralNetsweightMatrix_24_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_24_3 = io_inConf_bits_confneuralNetsweightMatrix_24_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_25_0 = io_inConf_bits_confneuralNetsweightMatrix_25_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_25_1 = io_inConf_bits_confneuralNetsweightMatrix_25_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_25_2 = io_inConf_bits_confneuralNetsweightMatrix_25_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_25_3 = io_inConf_bits_confneuralNetsweightMatrix_25_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_26_0 = io_inConf_bits_confneuralNetsweightMatrix_26_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_26_1 = io_inConf_bits_confneuralNetsweightMatrix_26_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_26_2 = io_inConf_bits_confneuralNetsweightMatrix_26_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_26_3 = io_inConf_bits_confneuralNetsweightMatrix_26_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_27_0 = io_inConf_bits_confneuralNetsweightMatrix_27_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_27_1 = io_inConf_bits_confneuralNetsweightMatrix_27_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_27_2 = io_inConf_bits_confneuralNetsweightMatrix_27_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_27_3 = io_inConf_bits_confneuralNetsweightMatrix_27_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_28_0 = io_inConf_bits_confneuralNetsweightMatrix_28_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_28_1 = io_inConf_bits_confneuralNetsweightMatrix_28_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_28_2 = io_inConf_bits_confneuralNetsweightMatrix_28_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_28_3 = io_inConf_bits_confneuralNetsweightMatrix_28_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_29_0 = io_inConf_bits_confneuralNetsweightMatrix_29_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_29_1 = io_inConf_bits_confneuralNetsweightMatrix_29_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_29_2 = io_inConf_bits_confneuralNetsweightMatrix_29_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_29_3 = io_inConf_bits_confneuralNetsweightMatrix_29_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_30_0 = io_inConf_bits_confneuralNetsweightMatrix_30_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_30_1 = io_inConf_bits_confneuralNetsweightMatrix_30_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_30_2 = io_inConf_bits_confneuralNetsweightMatrix_30_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_30_3 = io_inConf_bits_confneuralNetsweightMatrix_30_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_31_0 = io_inConf_bits_confneuralNetsweightMatrix_31_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_31_1 = io_inConf_bits_confneuralNetsweightMatrix_31_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_31_2 = io_inConf_bits_confneuralNetsweightMatrix_31_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_31_3 = io_inConf_bits_confneuralNetsweightMatrix_31_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_32_0 = io_inConf_bits_confneuralNetsweightMatrix_32_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_32_1 = io_inConf_bits_confneuralNetsweightMatrix_32_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_32_2 = io_inConf_bits_confneuralNetsweightMatrix_32_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_32_3 = io_inConf_bits_confneuralNetsweightMatrix_32_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_33_0 = io_inConf_bits_confneuralNetsweightMatrix_33_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_33_1 = io_inConf_bits_confneuralNetsweightMatrix_33_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_33_2 = io_inConf_bits_confneuralNetsweightMatrix_33_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_33_3 = io_inConf_bits_confneuralNetsweightMatrix_33_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_34_0 = io_inConf_bits_confneuralNetsweightMatrix_34_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_34_1 = io_inConf_bits_confneuralNetsweightMatrix_34_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_34_2 = io_inConf_bits_confneuralNetsweightMatrix_34_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_34_3 = io_inConf_bits_confneuralNetsweightMatrix_34_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_35_0 = io_inConf_bits_confneuralNetsweightMatrix_35_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_35_1 = io_inConf_bits_confneuralNetsweightMatrix_35_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_35_2 = io_inConf_bits_confneuralNetsweightMatrix_35_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_35_3 = io_inConf_bits_confneuralNetsweightMatrix_35_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_36_0 = io_inConf_bits_confneuralNetsweightMatrix_36_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_36_1 = io_inConf_bits_confneuralNetsweightMatrix_36_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_36_2 = io_inConf_bits_confneuralNetsweightMatrix_36_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_36_3 = io_inConf_bits_confneuralNetsweightMatrix_36_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_37_0 = io_inConf_bits_confneuralNetsweightMatrix_37_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_37_1 = io_inConf_bits_confneuralNetsweightMatrix_37_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_37_2 = io_inConf_bits_confneuralNetsweightMatrix_37_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_37_3 = io_inConf_bits_confneuralNetsweightMatrix_37_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_38_0 = io_inConf_bits_confneuralNetsweightMatrix_38_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_38_1 = io_inConf_bits_confneuralNetsweightMatrix_38_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_38_2 = io_inConf_bits_confneuralNetsweightMatrix_38_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_38_3 = io_inConf_bits_confneuralNetsweightMatrix_38_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_39_0 = io_inConf_bits_confneuralNetsweightMatrix_39_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_39_1 = io_inConf_bits_confneuralNetsweightMatrix_39_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_39_2 = io_inConf_bits_confneuralNetsweightMatrix_39_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_39_3 = io_inConf_bits_confneuralNetsweightMatrix_39_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_40_0 = io_inConf_bits_confneuralNetsweightMatrix_40_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_40_1 = io_inConf_bits_confneuralNetsweightMatrix_40_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_40_2 = io_inConf_bits_confneuralNetsweightMatrix_40_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_40_3 = io_inConf_bits_confneuralNetsweightMatrix_40_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_41_0 = io_inConf_bits_confneuralNetsweightMatrix_41_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_41_1 = io_inConf_bits_confneuralNetsweightMatrix_41_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_41_2 = io_inConf_bits_confneuralNetsweightMatrix_41_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_41_3 = io_inConf_bits_confneuralNetsweightMatrix_41_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_42_0 = io_inConf_bits_confneuralNetsweightMatrix_42_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_42_1 = io_inConf_bits_confneuralNetsweightMatrix_42_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_42_2 = io_inConf_bits_confneuralNetsweightMatrix_42_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_42_3 = io_inConf_bits_confneuralNetsweightMatrix_42_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_43_0 = io_inConf_bits_confneuralNetsweightMatrix_43_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_43_1 = io_inConf_bits_confneuralNetsweightMatrix_43_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_43_2 = io_inConf_bits_confneuralNetsweightMatrix_43_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_43_3 = io_inConf_bits_confneuralNetsweightMatrix_43_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_44_0 = io_inConf_bits_confneuralNetsweightMatrix_44_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_44_1 = io_inConf_bits_confneuralNetsweightMatrix_44_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_44_2 = io_inConf_bits_confneuralNetsweightMatrix_44_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_44_3 = io_inConf_bits_confneuralNetsweightMatrix_44_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_45_0 = io_inConf_bits_confneuralNetsweightMatrix_45_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_45_1 = io_inConf_bits_confneuralNetsweightMatrix_45_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_45_2 = io_inConf_bits_confneuralNetsweightMatrix_45_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_45_3 = io_inConf_bits_confneuralNetsweightMatrix_45_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_46_0 = io_inConf_bits_confneuralNetsweightMatrix_46_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_46_1 = io_inConf_bits_confneuralNetsweightMatrix_46_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_46_2 = io_inConf_bits_confneuralNetsweightMatrix_46_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_46_3 = io_inConf_bits_confneuralNetsweightMatrix_46_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_47_0 = io_inConf_bits_confneuralNetsweightMatrix_47_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_47_1 = io_inConf_bits_confneuralNetsweightMatrix_47_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_47_2 = io_inConf_bits_confneuralNetsweightMatrix_47_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_47_3 = io_inConf_bits_confneuralNetsweightMatrix_47_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_48_0 = io_inConf_bits_confneuralNetsweightMatrix_48_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_48_1 = io_inConf_bits_confneuralNetsweightMatrix_48_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_48_2 = io_inConf_bits_confneuralNetsweightMatrix_48_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_48_3 = io_inConf_bits_confneuralNetsweightMatrix_48_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_49_0 = io_inConf_bits_confneuralNetsweightMatrix_49_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_49_1 = io_inConf_bits_confneuralNetsweightMatrix_49_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_49_2 = io_inConf_bits_confneuralNetsweightMatrix_49_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_49_3 = io_inConf_bits_confneuralNetsweightMatrix_49_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_50_0 = io_inConf_bits_confneuralNetsweightMatrix_50_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_50_1 = io_inConf_bits_confneuralNetsweightMatrix_50_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_50_2 = io_inConf_bits_confneuralNetsweightMatrix_50_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_50_3 = io_inConf_bits_confneuralNetsweightMatrix_50_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_51_0 = io_inConf_bits_confneuralNetsweightMatrix_51_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_51_1 = io_inConf_bits_confneuralNetsweightMatrix_51_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_51_2 = io_inConf_bits_confneuralNetsweightMatrix_51_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_51_3 = io_inConf_bits_confneuralNetsweightMatrix_51_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_52_0 = io_inConf_bits_confneuralNetsweightMatrix_52_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_52_1 = io_inConf_bits_confneuralNetsweightMatrix_52_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_52_2 = io_inConf_bits_confneuralNetsweightMatrix_52_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_52_3 = io_inConf_bits_confneuralNetsweightMatrix_52_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_53_0 = io_inConf_bits_confneuralNetsweightMatrix_53_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_53_1 = io_inConf_bits_confneuralNetsweightMatrix_53_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_53_2 = io_inConf_bits_confneuralNetsweightMatrix_53_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_53_3 = io_inConf_bits_confneuralNetsweightMatrix_53_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_54_0 = io_inConf_bits_confneuralNetsweightMatrix_54_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_54_1 = io_inConf_bits_confneuralNetsweightMatrix_54_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_54_2 = io_inConf_bits_confneuralNetsweightMatrix_54_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_54_3 = io_inConf_bits_confneuralNetsweightMatrix_54_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_55_0 = io_inConf_bits_confneuralNetsweightMatrix_55_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_55_1 = io_inConf_bits_confneuralNetsweightMatrix_55_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_55_2 = io_inConf_bits_confneuralNetsweightMatrix_55_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_55_3 = io_inConf_bits_confneuralNetsweightMatrix_55_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_56_0 = io_inConf_bits_confneuralNetsweightMatrix_56_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_56_1 = io_inConf_bits_confneuralNetsweightMatrix_56_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_56_2 = io_inConf_bits_confneuralNetsweightMatrix_56_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_56_3 = io_inConf_bits_confneuralNetsweightMatrix_56_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_57_0 = io_inConf_bits_confneuralNetsweightMatrix_57_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_57_1 = io_inConf_bits_confneuralNetsweightMatrix_57_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_57_2 = io_inConf_bits_confneuralNetsweightMatrix_57_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_57_3 = io_inConf_bits_confneuralNetsweightMatrix_57_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_58_0 = io_inConf_bits_confneuralNetsweightMatrix_58_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_58_1 = io_inConf_bits_confneuralNetsweightMatrix_58_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_58_2 = io_inConf_bits_confneuralNetsweightMatrix_58_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_58_3 = io_inConf_bits_confneuralNetsweightMatrix_58_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_59_0 = io_inConf_bits_confneuralNetsweightMatrix_59_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_59_1 = io_inConf_bits_confneuralNetsweightMatrix_59_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_59_2 = io_inConf_bits_confneuralNetsweightMatrix_59_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_59_3 = io_inConf_bits_confneuralNetsweightMatrix_59_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_60_0 = io_inConf_bits_confneuralNetsweightMatrix_60_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_60_1 = io_inConf_bits_confneuralNetsweightMatrix_60_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_60_2 = io_inConf_bits_confneuralNetsweightMatrix_60_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_60_3 = io_inConf_bits_confneuralNetsweightMatrix_60_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_61_0 = io_inConf_bits_confneuralNetsweightMatrix_61_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_61_1 = io_inConf_bits_confneuralNetsweightMatrix_61_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_61_2 = io_inConf_bits_confneuralNetsweightMatrix_61_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_61_3 = io_inConf_bits_confneuralNetsweightMatrix_61_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_62_0 = io_inConf_bits_confneuralNetsweightMatrix_62_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_62_1 = io_inConf_bits_confneuralNetsweightMatrix_62_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_62_2 = io_inConf_bits_confneuralNetsweightMatrix_62_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_62_3 = io_inConf_bits_confneuralNetsweightMatrix_62_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_63_0 = io_inConf_bits_confneuralNetsweightMatrix_63_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_63_1 = io_inConf_bits_confneuralNetsweightMatrix_63_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_63_2 = io_inConf_bits_confneuralNetsweightMatrix_63_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_63_3 = io_inConf_bits_confneuralNetsweightMatrix_63_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_64_0 = io_inConf_bits_confneuralNetsweightMatrix_64_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_64_1 = io_inConf_bits_confneuralNetsweightMatrix_64_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_64_2 = io_inConf_bits_confneuralNetsweightMatrix_64_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_64_3 = io_inConf_bits_confneuralNetsweightMatrix_64_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_65_0 = io_inConf_bits_confneuralNetsweightMatrix_65_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_65_1 = io_inConf_bits_confneuralNetsweightMatrix_65_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_65_2 = io_inConf_bits_confneuralNetsweightMatrix_65_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_65_3 = io_inConf_bits_confneuralNetsweightMatrix_65_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_66_0 = io_inConf_bits_confneuralNetsweightMatrix_66_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_66_1 = io_inConf_bits_confneuralNetsweightMatrix_66_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_66_2 = io_inConf_bits_confneuralNetsweightMatrix_66_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_66_3 = io_inConf_bits_confneuralNetsweightMatrix_66_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_67_0 = io_inConf_bits_confneuralNetsweightMatrix_67_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_67_1 = io_inConf_bits_confneuralNetsweightMatrix_67_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_67_2 = io_inConf_bits_confneuralNetsweightMatrix_67_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_67_3 = io_inConf_bits_confneuralNetsweightMatrix_67_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_68_0 = io_inConf_bits_confneuralNetsweightMatrix_68_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_68_1 = io_inConf_bits_confneuralNetsweightMatrix_68_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_68_2 = io_inConf_bits_confneuralNetsweightMatrix_68_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_68_3 = io_inConf_bits_confneuralNetsweightMatrix_68_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_69_0 = io_inConf_bits_confneuralNetsweightMatrix_69_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_69_1 = io_inConf_bits_confneuralNetsweightMatrix_69_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_69_2 = io_inConf_bits_confneuralNetsweightMatrix_69_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_69_3 = io_inConf_bits_confneuralNetsweightMatrix_69_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_70_0 = io_inConf_bits_confneuralNetsweightMatrix_70_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_70_1 = io_inConf_bits_confneuralNetsweightMatrix_70_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_70_2 = io_inConf_bits_confneuralNetsweightMatrix_70_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_70_3 = io_inConf_bits_confneuralNetsweightMatrix_70_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_71_0 = io_inConf_bits_confneuralNetsweightMatrix_71_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_71_1 = io_inConf_bits_confneuralNetsweightMatrix_71_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_71_2 = io_inConf_bits_confneuralNetsweightMatrix_71_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_71_3 = io_inConf_bits_confneuralNetsweightMatrix_71_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_72_0 = io_inConf_bits_confneuralNetsweightMatrix_72_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_72_1 = io_inConf_bits_confneuralNetsweightMatrix_72_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_72_2 = io_inConf_bits_confneuralNetsweightMatrix_72_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_72_3 = io_inConf_bits_confneuralNetsweightMatrix_72_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_73_0 = io_inConf_bits_confneuralNetsweightMatrix_73_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_73_1 = io_inConf_bits_confneuralNetsweightMatrix_73_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_73_2 = io_inConf_bits_confneuralNetsweightMatrix_73_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_73_3 = io_inConf_bits_confneuralNetsweightMatrix_73_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_74_0 = io_inConf_bits_confneuralNetsweightMatrix_74_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_74_1 = io_inConf_bits_confneuralNetsweightMatrix_74_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_74_2 = io_inConf_bits_confneuralNetsweightMatrix_74_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_74_3 = io_inConf_bits_confneuralNetsweightMatrix_74_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_75_0 = io_inConf_bits_confneuralNetsweightMatrix_75_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_75_1 = io_inConf_bits_confneuralNetsweightMatrix_75_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_75_2 = io_inConf_bits_confneuralNetsweightMatrix_75_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_75_3 = io_inConf_bits_confneuralNetsweightMatrix_75_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_76_0 = io_inConf_bits_confneuralNetsweightMatrix_76_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_76_1 = io_inConf_bits_confneuralNetsweightMatrix_76_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_76_2 = io_inConf_bits_confneuralNetsweightMatrix_76_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_76_3 = io_inConf_bits_confneuralNetsweightMatrix_76_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_77_0 = io_inConf_bits_confneuralNetsweightMatrix_77_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_77_1 = io_inConf_bits_confneuralNetsweightMatrix_77_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_77_2 = io_inConf_bits_confneuralNetsweightMatrix_77_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_77_3 = io_inConf_bits_confneuralNetsweightMatrix_77_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_78_0 = io_inConf_bits_confneuralNetsweightMatrix_78_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_78_1 = io_inConf_bits_confneuralNetsweightMatrix_78_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_78_2 = io_inConf_bits_confneuralNetsweightMatrix_78_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_78_3 = io_inConf_bits_confneuralNetsweightMatrix_78_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_79_0 = io_inConf_bits_confneuralNetsweightMatrix_79_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_79_1 = io_inConf_bits_confneuralNetsweightMatrix_79_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_79_2 = io_inConf_bits_confneuralNetsweightMatrix_79_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_79_3 = io_inConf_bits_confneuralNetsweightMatrix_79_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_80_0 = io_inConf_bits_confneuralNetsweightMatrix_80_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_80_1 = io_inConf_bits_confneuralNetsweightMatrix_80_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_80_2 = io_inConf_bits_confneuralNetsweightMatrix_80_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_80_3 = io_inConf_bits_confneuralNetsweightMatrix_80_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_81_0 = io_inConf_bits_confneuralNetsweightMatrix_81_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_81_1 = io_inConf_bits_confneuralNetsweightMatrix_81_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_81_2 = io_inConf_bits_confneuralNetsweightMatrix_81_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_81_3 = io_inConf_bits_confneuralNetsweightMatrix_81_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_82_0 = io_inConf_bits_confneuralNetsweightMatrix_82_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_82_1 = io_inConf_bits_confneuralNetsweightMatrix_82_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_82_2 = io_inConf_bits_confneuralNetsweightMatrix_82_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_82_3 = io_inConf_bits_confneuralNetsweightMatrix_82_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_83_0 = io_inConf_bits_confneuralNetsweightMatrix_83_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_83_1 = io_inConf_bits_confneuralNetsweightMatrix_83_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_83_2 = io_inConf_bits_confneuralNetsweightMatrix_83_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_83_3 = io_inConf_bits_confneuralNetsweightMatrix_83_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_84_0 = io_inConf_bits_confneuralNetsweightMatrix_84_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_84_1 = io_inConf_bits_confneuralNetsweightMatrix_84_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_84_2 = io_inConf_bits_confneuralNetsweightMatrix_84_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_84_3 = io_inConf_bits_confneuralNetsweightMatrix_84_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_85_0 = io_inConf_bits_confneuralNetsweightMatrix_85_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_85_1 = io_inConf_bits_confneuralNetsweightMatrix_85_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_85_2 = io_inConf_bits_confneuralNetsweightMatrix_85_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_85_3 = io_inConf_bits_confneuralNetsweightMatrix_85_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_86_0 = io_inConf_bits_confneuralNetsweightMatrix_86_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_86_1 = io_inConf_bits_confneuralNetsweightMatrix_86_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_86_2 = io_inConf_bits_confneuralNetsweightMatrix_86_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_86_3 = io_inConf_bits_confneuralNetsweightMatrix_86_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_87_0 = io_inConf_bits_confneuralNetsweightMatrix_87_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_87_1 = io_inConf_bits_confneuralNetsweightMatrix_87_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_87_2 = io_inConf_bits_confneuralNetsweightMatrix_87_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_87_3 = io_inConf_bits_confneuralNetsweightMatrix_87_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_88_0 = io_inConf_bits_confneuralNetsweightMatrix_88_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_88_1 = io_inConf_bits_confneuralNetsweightMatrix_88_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_88_2 = io_inConf_bits_confneuralNetsweightMatrix_88_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_88_3 = io_inConf_bits_confneuralNetsweightMatrix_88_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_89_0 = io_inConf_bits_confneuralNetsweightMatrix_89_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_89_1 = io_inConf_bits_confneuralNetsweightMatrix_89_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_89_2 = io_inConf_bits_confneuralNetsweightMatrix_89_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_89_3 = io_inConf_bits_confneuralNetsweightMatrix_89_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_90_0 = io_inConf_bits_confneuralNetsweightMatrix_90_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_90_1 = io_inConf_bits_confneuralNetsweightMatrix_90_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_90_2 = io_inConf_bits_confneuralNetsweightMatrix_90_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_90_3 = io_inConf_bits_confneuralNetsweightMatrix_90_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_91_0 = io_inConf_bits_confneuralNetsweightMatrix_91_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_91_1 = io_inConf_bits_confneuralNetsweightMatrix_91_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_91_2 = io_inConf_bits_confneuralNetsweightMatrix_91_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_91_3 = io_inConf_bits_confneuralNetsweightMatrix_91_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_92_0 = io_inConf_bits_confneuralNetsweightMatrix_92_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_92_1 = io_inConf_bits_confneuralNetsweightMatrix_92_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_92_2 = io_inConf_bits_confneuralNetsweightMatrix_92_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_92_3 = io_inConf_bits_confneuralNetsweightMatrix_92_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_93_0 = io_inConf_bits_confneuralNetsweightMatrix_93_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_93_1 = io_inConf_bits_confneuralNetsweightMatrix_93_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_93_2 = io_inConf_bits_confneuralNetsweightMatrix_93_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_93_3 = io_inConf_bits_confneuralNetsweightMatrix_93_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_94_0 = io_inConf_bits_confneuralNetsweightMatrix_94_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_94_1 = io_inConf_bits_confneuralNetsweightMatrix_94_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_94_2 = io_inConf_bits_confneuralNetsweightMatrix_94_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_94_3 = io_inConf_bits_confneuralNetsweightMatrix_94_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_95_0 = io_inConf_bits_confneuralNetsweightMatrix_95_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_95_1 = io_inConf_bits_confneuralNetsweightMatrix_95_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_95_2 = io_inConf_bits_confneuralNetsweightMatrix_95_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_95_3 = io_inConf_bits_confneuralNetsweightMatrix_95_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_96_0 = io_inConf_bits_confneuralNetsweightMatrix_96_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_96_1 = io_inConf_bits_confneuralNetsweightMatrix_96_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_96_2 = io_inConf_bits_confneuralNetsweightMatrix_96_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_96_3 = io_inConf_bits_confneuralNetsweightMatrix_96_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_97_0 = io_inConf_bits_confneuralNetsweightMatrix_97_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_97_1 = io_inConf_bits_confneuralNetsweightMatrix_97_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_97_2 = io_inConf_bits_confneuralNetsweightMatrix_97_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_97_3 = io_inConf_bits_confneuralNetsweightMatrix_97_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_98_0 = io_inConf_bits_confneuralNetsweightMatrix_98_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_98_1 = io_inConf_bits_confneuralNetsweightMatrix_98_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_98_2 = io_inConf_bits_confneuralNetsweightMatrix_98_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_98_3 = io_inConf_bits_confneuralNetsweightMatrix_98_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_99_0 = io_inConf_bits_confneuralNetsweightMatrix_99_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_99_1 = io_inConf_bits_confneuralNetsweightMatrix_99_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_99_2 = io_inConf_bits_confneuralNetsweightMatrix_99_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightMatrix_99_3 = io_inConf_bits_confneuralNetsweightMatrix_99_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_weightVec_0 = io_inConf_bits_confneuralNetsweightVec_0; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_1 = io_inConf_bits_confneuralNetsweightVec_1; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_2 = io_inConf_bits_confneuralNetsweightVec_2; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_3 = io_inConf_bits_confneuralNetsweightVec_3; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_4 = io_inConf_bits_confneuralNetsweightVec_4; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_5 = io_inConf_bits_confneuralNetsweightVec_5; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_6 = io_inConf_bits_confneuralNetsweightVec_6; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_7 = io_inConf_bits_confneuralNetsweightVec_7; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_8 = io_inConf_bits_confneuralNetsweightVec_8; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_9 = io_inConf_bits_confneuralNetsweightVec_9; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_10 = io_inConf_bits_confneuralNetsweightVec_10; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_11 = io_inConf_bits_confneuralNetsweightVec_11; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_12 = io_inConf_bits_confneuralNetsweightVec_12; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_13 = io_inConf_bits_confneuralNetsweightVec_13; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_14 = io_inConf_bits_confneuralNetsweightVec_14; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_15 = io_inConf_bits_confneuralNetsweightVec_15; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_16 = io_inConf_bits_confneuralNetsweightVec_16; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_17 = io_inConf_bits_confneuralNetsweightVec_17; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_18 = io_inConf_bits_confneuralNetsweightVec_18; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_19 = io_inConf_bits_confneuralNetsweightVec_19; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_20 = io_inConf_bits_confneuralNetsweightVec_20; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_21 = io_inConf_bits_confneuralNetsweightVec_21; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_22 = io_inConf_bits_confneuralNetsweightVec_22; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_23 = io_inConf_bits_confneuralNetsweightVec_23; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_24 = io_inConf_bits_confneuralNetsweightVec_24; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_25 = io_inConf_bits_confneuralNetsweightVec_25; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_26 = io_inConf_bits_confneuralNetsweightVec_26; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_27 = io_inConf_bits_confneuralNetsweightVec_27; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_28 = io_inConf_bits_confneuralNetsweightVec_28; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_29 = io_inConf_bits_confneuralNetsweightVec_29; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_30 = io_inConf_bits_confneuralNetsweightVec_30; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_31 = io_inConf_bits_confneuralNetsweightVec_31; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_32 = io_inConf_bits_confneuralNetsweightVec_32; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_33 = io_inConf_bits_confneuralNetsweightVec_33; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_34 = io_inConf_bits_confneuralNetsweightVec_34; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_35 = io_inConf_bits_confneuralNetsweightVec_35; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_36 = io_inConf_bits_confneuralNetsweightVec_36; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_37 = io_inConf_bits_confneuralNetsweightVec_37; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_38 = io_inConf_bits_confneuralNetsweightVec_38; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_39 = io_inConf_bits_confneuralNetsweightVec_39; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_40 = io_inConf_bits_confneuralNetsweightVec_40; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_41 = io_inConf_bits_confneuralNetsweightVec_41; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_42 = io_inConf_bits_confneuralNetsweightVec_42; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_43 = io_inConf_bits_confneuralNetsweightVec_43; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_44 = io_inConf_bits_confneuralNetsweightVec_44; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_45 = io_inConf_bits_confneuralNetsweightVec_45; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_46 = io_inConf_bits_confneuralNetsweightVec_46; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_47 = io_inConf_bits_confneuralNetsweightVec_47; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_48 = io_inConf_bits_confneuralNetsweightVec_48; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_49 = io_inConf_bits_confneuralNetsweightVec_49; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_50 = io_inConf_bits_confneuralNetsweightVec_50; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_51 = io_inConf_bits_confneuralNetsweightVec_51; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_52 = io_inConf_bits_confneuralNetsweightVec_52; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_53 = io_inConf_bits_confneuralNetsweightVec_53; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_54 = io_inConf_bits_confneuralNetsweightVec_54; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_55 = io_inConf_bits_confneuralNetsweightVec_55; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_56 = io_inConf_bits_confneuralNetsweightVec_56; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_57 = io_inConf_bits_confneuralNetsweightVec_57; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_58 = io_inConf_bits_confneuralNetsweightVec_58; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_59 = io_inConf_bits_confneuralNetsweightVec_59; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_60 = io_inConf_bits_confneuralNetsweightVec_60; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_61 = io_inConf_bits_confneuralNetsweightVec_61; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_62 = io_inConf_bits_confneuralNetsweightVec_62; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_63 = io_inConf_bits_confneuralNetsweightVec_63; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_64 = io_inConf_bits_confneuralNetsweightVec_64; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_65 = io_inConf_bits_confneuralNetsweightVec_65; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_66 = io_inConf_bits_confneuralNetsweightVec_66; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_67 = io_inConf_bits_confneuralNetsweightVec_67; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_68 = io_inConf_bits_confneuralNetsweightVec_68; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_69 = io_inConf_bits_confneuralNetsweightVec_69; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_70 = io_inConf_bits_confneuralNetsweightVec_70; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_71 = io_inConf_bits_confneuralNetsweightVec_71; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_72 = io_inConf_bits_confneuralNetsweightVec_72; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_73 = io_inConf_bits_confneuralNetsweightVec_73; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_74 = io_inConf_bits_confneuralNetsweightVec_74; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_75 = io_inConf_bits_confneuralNetsweightVec_75; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_76 = io_inConf_bits_confneuralNetsweightVec_76; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_77 = io_inConf_bits_confneuralNetsweightVec_77; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_78 = io_inConf_bits_confneuralNetsweightVec_78; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_79 = io_inConf_bits_confneuralNetsweightVec_79; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_80 = io_inConf_bits_confneuralNetsweightVec_80; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_81 = io_inConf_bits_confneuralNetsweightVec_81; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_82 = io_inConf_bits_confneuralNetsweightVec_82; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_83 = io_inConf_bits_confneuralNetsweightVec_83; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_84 = io_inConf_bits_confneuralNetsweightVec_84; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_85 = io_inConf_bits_confneuralNetsweightVec_85; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_86 = io_inConf_bits_confneuralNetsweightVec_86; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_87 = io_inConf_bits_confneuralNetsweightVec_87; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_88 = io_inConf_bits_confneuralNetsweightVec_88; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_89 = io_inConf_bits_confneuralNetsweightVec_89; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_90 = io_inConf_bits_confneuralNetsweightVec_90; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_91 = io_inConf_bits_confneuralNetsweightVec_91; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_92 = io_inConf_bits_confneuralNetsweightVec_92; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_93 = io_inConf_bits_confneuralNetsweightVec_93; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_94 = io_inConf_bits_confneuralNetsweightVec_94; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_95 = io_inConf_bits_confneuralNetsweightVec_95; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_96 = io_inConf_bits_confneuralNetsweightVec_96; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_97 = io_inConf_bits_confneuralNetsweightVec_97; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_98 = io_inConf_bits_confneuralNetsweightVec_98; // @[Wellness.scala 337:27]
  assign neuralNets_io_weightVec_99 = io_inConf_bits_confneuralNetsweightVec_99; // @[Wellness.scala 337:27]
  assign neuralNets_io_biasVec_0 = io_inConf_bits_confneuralNetsbiasVec_0; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_1 = io_inConf_bits_confneuralNetsbiasVec_1; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_2 = io_inConf_bits_confneuralNetsbiasVec_2; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_3 = io_inConf_bits_confneuralNetsbiasVec_3; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_4 = io_inConf_bits_confneuralNetsbiasVec_4; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_5 = io_inConf_bits_confneuralNetsbiasVec_5; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_6 = io_inConf_bits_confneuralNetsbiasVec_6; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_7 = io_inConf_bits_confneuralNetsbiasVec_7; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_8 = io_inConf_bits_confneuralNetsbiasVec_8; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_9 = io_inConf_bits_confneuralNetsbiasVec_9; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_10 = io_inConf_bits_confneuralNetsbiasVec_10; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_11 = io_inConf_bits_confneuralNetsbiasVec_11; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_12 = io_inConf_bits_confneuralNetsbiasVec_12; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_13 = io_inConf_bits_confneuralNetsbiasVec_13; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_14 = io_inConf_bits_confneuralNetsbiasVec_14; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_15 = io_inConf_bits_confneuralNetsbiasVec_15; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_16 = io_inConf_bits_confneuralNetsbiasVec_16; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_17 = io_inConf_bits_confneuralNetsbiasVec_17; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_18 = io_inConf_bits_confneuralNetsbiasVec_18; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_19 = io_inConf_bits_confneuralNetsbiasVec_19; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_20 = io_inConf_bits_confneuralNetsbiasVec_20; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_21 = io_inConf_bits_confneuralNetsbiasVec_21; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_22 = io_inConf_bits_confneuralNetsbiasVec_22; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_23 = io_inConf_bits_confneuralNetsbiasVec_23; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_24 = io_inConf_bits_confneuralNetsbiasVec_24; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_25 = io_inConf_bits_confneuralNetsbiasVec_25; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_26 = io_inConf_bits_confneuralNetsbiasVec_26; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_27 = io_inConf_bits_confneuralNetsbiasVec_27; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_28 = io_inConf_bits_confneuralNetsbiasVec_28; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_29 = io_inConf_bits_confneuralNetsbiasVec_29; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_30 = io_inConf_bits_confneuralNetsbiasVec_30; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_31 = io_inConf_bits_confneuralNetsbiasVec_31; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_32 = io_inConf_bits_confneuralNetsbiasVec_32; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_33 = io_inConf_bits_confneuralNetsbiasVec_33; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_34 = io_inConf_bits_confneuralNetsbiasVec_34; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_35 = io_inConf_bits_confneuralNetsbiasVec_35; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_36 = io_inConf_bits_confneuralNetsbiasVec_36; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_37 = io_inConf_bits_confneuralNetsbiasVec_37; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_38 = io_inConf_bits_confneuralNetsbiasVec_38; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_39 = io_inConf_bits_confneuralNetsbiasVec_39; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_40 = io_inConf_bits_confneuralNetsbiasVec_40; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_41 = io_inConf_bits_confneuralNetsbiasVec_41; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_42 = io_inConf_bits_confneuralNetsbiasVec_42; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_43 = io_inConf_bits_confneuralNetsbiasVec_43; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_44 = io_inConf_bits_confneuralNetsbiasVec_44; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_45 = io_inConf_bits_confneuralNetsbiasVec_45; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_46 = io_inConf_bits_confneuralNetsbiasVec_46; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_47 = io_inConf_bits_confneuralNetsbiasVec_47; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_48 = io_inConf_bits_confneuralNetsbiasVec_48; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_49 = io_inConf_bits_confneuralNetsbiasVec_49; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_50 = io_inConf_bits_confneuralNetsbiasVec_50; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_51 = io_inConf_bits_confneuralNetsbiasVec_51; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_52 = io_inConf_bits_confneuralNetsbiasVec_52; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_53 = io_inConf_bits_confneuralNetsbiasVec_53; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_54 = io_inConf_bits_confneuralNetsbiasVec_54; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_55 = io_inConf_bits_confneuralNetsbiasVec_55; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_56 = io_inConf_bits_confneuralNetsbiasVec_56; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_57 = io_inConf_bits_confneuralNetsbiasVec_57; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_58 = io_inConf_bits_confneuralNetsbiasVec_58; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_59 = io_inConf_bits_confneuralNetsbiasVec_59; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_60 = io_inConf_bits_confneuralNetsbiasVec_60; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_61 = io_inConf_bits_confneuralNetsbiasVec_61; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_62 = io_inConf_bits_confneuralNetsbiasVec_62; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_63 = io_inConf_bits_confneuralNetsbiasVec_63; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_64 = io_inConf_bits_confneuralNetsbiasVec_64; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_65 = io_inConf_bits_confneuralNetsbiasVec_65; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_66 = io_inConf_bits_confneuralNetsbiasVec_66; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_67 = io_inConf_bits_confneuralNetsbiasVec_67; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_68 = io_inConf_bits_confneuralNetsbiasVec_68; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_69 = io_inConf_bits_confneuralNetsbiasVec_69; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_70 = io_inConf_bits_confneuralNetsbiasVec_70; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_71 = io_inConf_bits_confneuralNetsbiasVec_71; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_72 = io_inConf_bits_confneuralNetsbiasVec_72; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_73 = io_inConf_bits_confneuralNetsbiasVec_73; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_74 = io_inConf_bits_confneuralNetsbiasVec_74; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_75 = io_inConf_bits_confneuralNetsbiasVec_75; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_76 = io_inConf_bits_confneuralNetsbiasVec_76; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_77 = io_inConf_bits_confneuralNetsbiasVec_77; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_78 = io_inConf_bits_confneuralNetsbiasVec_78; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_79 = io_inConf_bits_confneuralNetsbiasVec_79; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_80 = io_inConf_bits_confneuralNetsbiasVec_80; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_81 = io_inConf_bits_confneuralNetsbiasVec_81; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_82 = io_inConf_bits_confneuralNetsbiasVec_82; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_83 = io_inConf_bits_confneuralNetsbiasVec_83; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_84 = io_inConf_bits_confneuralNetsbiasVec_84; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_85 = io_inConf_bits_confneuralNetsbiasVec_85; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_86 = io_inConf_bits_confneuralNetsbiasVec_86; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_87 = io_inConf_bits_confneuralNetsbiasVec_87; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_88 = io_inConf_bits_confneuralNetsbiasVec_88; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_89 = io_inConf_bits_confneuralNetsbiasVec_89; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_90 = io_inConf_bits_confneuralNetsbiasVec_90; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_91 = io_inConf_bits_confneuralNetsbiasVec_91; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_92 = io_inConf_bits_confneuralNetsbiasVec_92; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_93 = io_inConf_bits_confneuralNetsbiasVec_93; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_94 = io_inConf_bits_confneuralNetsbiasVec_94; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_95 = io_inConf_bits_confneuralNetsbiasVec_95; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_96 = io_inConf_bits_confneuralNetsbiasVec_96; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_97 = io_inConf_bits_confneuralNetsbiasVec_97; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_98 = io_inConf_bits_confneuralNetsbiasVec_98; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasVec_99 = io_inConf_bits_confneuralNetsbiasVec_99; // @[Wellness.scala 338:25]
  assign neuralNets_io_biasScalar = io_inConf_bits_confneuralNetsbiasScalar_0; // @[Wellness.scala 339:28]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  lineLength1Reg1 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  lineLength1Valid1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    lineLength1Reg1 <= $signed(_T_22);
    lineLength1Valid1 <= lineLength1_io_out_valid;
  end
endmodule
module MemoryBuffer(
  input         clock,
  input         reset,
  input         io_in_valid,
  input  [31:0] io_in_bits,
  output [31:0] io_out_bits_0_0,
  output [31:0] io_out_bits_0_1,
  output [31:0] io_out_bits_0_2,
  output [31:0] io_out_bits_0_3,
  output [31:0] io_out_bits_1_0,
  output [31:0] io_out_bits_1_1,
  output [31:0] io_out_bits_1_2,
  output [31:0] io_out_bits_1_3,
  output [31:0] io_out_bits_2_0,
  output [31:0] io_out_bits_2_1,
  output [31:0] io_out_bits_2_2,
  output [31:0] io_out_bits_2_3,
  output [31:0] io_out_bits_3_0,
  output [31:0] io_out_bits_3_1,
  output [31:0] io_out_bits_3_2,
  output [31:0] io_out_bits_3_3,
  output [31:0] io_out_bits_4_0,
  output [31:0] io_out_bits_4_1,
  output [31:0] io_out_bits_4_2,
  output [31:0] io_out_bits_4_3,
  output [31:0] io_out_bits_5_0,
  output [31:0] io_out_bits_5_1,
  output [31:0] io_out_bits_5_2,
  output [31:0] io_out_bits_5_3,
  output [31:0] io_out_bits_6_0,
  output [31:0] io_out_bits_6_1,
  output [31:0] io_out_bits_6_2,
  output [31:0] io_out_bits_6_3,
  output [31:0] io_out_bits_7_0,
  output [31:0] io_out_bits_7_1,
  output [31:0] io_out_bits_7_2,
  output [31:0] io_out_bits_7_3,
  output [31:0] io_out_bits_8_0,
  output [31:0] io_out_bits_8_1,
  output [31:0] io_out_bits_8_2,
  output [31:0] io_out_bits_8_3,
  output [31:0] io_out_bits_9_0,
  output [31:0] io_out_bits_9_1,
  output [31:0] io_out_bits_9_2,
  output [31:0] io_out_bits_9_3,
  output [31:0] io_out_bits_10_0,
  output [31:0] io_out_bits_10_1,
  output [31:0] io_out_bits_10_2,
  output [31:0] io_out_bits_10_3,
  output [31:0] io_out_bits_11_0,
  output [31:0] io_out_bits_11_1,
  output [31:0] io_out_bits_11_2,
  output [31:0] io_out_bits_11_3,
  output [31:0] io_out_bits_12_0,
  output [31:0] io_out_bits_12_1,
  output [31:0] io_out_bits_12_2,
  output [31:0] io_out_bits_12_3,
  output [31:0] io_out_bits_13_0,
  output [31:0] io_out_bits_13_1,
  output [31:0] io_out_bits_13_2,
  output [31:0] io_out_bits_13_3,
  output [31:0] io_out_bits_14_0,
  output [31:0] io_out_bits_14_1,
  output [31:0] io_out_bits_14_2,
  output [31:0] io_out_bits_14_3,
  output [31:0] io_out_bits_15_0,
  output [31:0] io_out_bits_15_1,
  output [31:0] io_out_bits_15_2,
  output [31:0] io_out_bits_15_3,
  output [31:0] io_out_bits_16_0,
  output [31:0] io_out_bits_16_1,
  output [31:0] io_out_bits_16_2,
  output [31:0] io_out_bits_16_3,
  output [31:0] io_out_bits_17_0,
  output [31:0] io_out_bits_17_1,
  output [31:0] io_out_bits_17_2,
  output [31:0] io_out_bits_17_3,
  output [31:0] io_out_bits_18_0,
  output [31:0] io_out_bits_18_1,
  output [31:0] io_out_bits_18_2,
  output [31:0] io_out_bits_18_3,
  output [31:0] io_out_bits_19_0,
  output [31:0] io_out_bits_19_1,
  output [31:0] io_out_bits_19_2,
  output [31:0] io_out_bits_19_3,
  output [31:0] io_out_bits_20_0,
  output [31:0] io_out_bits_20_1,
  output [31:0] io_out_bits_20_2,
  output [31:0] io_out_bits_20_3,
  output [31:0] io_out_bits_21_0,
  output [31:0] io_out_bits_21_1,
  output [31:0] io_out_bits_21_2,
  output [31:0] io_out_bits_21_3,
  output [31:0] io_out_bits_22_0,
  output [31:0] io_out_bits_22_1,
  output [31:0] io_out_bits_22_2,
  output [31:0] io_out_bits_22_3,
  output [31:0] io_out_bits_23_0,
  output [31:0] io_out_bits_23_1,
  output [31:0] io_out_bits_23_2,
  output [31:0] io_out_bits_23_3,
  output [31:0] io_out_bits_24_0,
  output [31:0] io_out_bits_24_1,
  output [31:0] io_out_bits_24_2,
  output [31:0] io_out_bits_24_3,
  output [31:0] io_out_bits_25_0,
  output [31:0] io_out_bits_25_1,
  output [31:0] io_out_bits_25_2,
  output [31:0] io_out_bits_25_3,
  output [31:0] io_out_bits_26_0,
  output [31:0] io_out_bits_26_1,
  output [31:0] io_out_bits_26_2,
  output [31:0] io_out_bits_26_3,
  output [31:0] io_out_bits_27_0,
  output [31:0] io_out_bits_27_1,
  output [31:0] io_out_bits_27_2,
  output [31:0] io_out_bits_27_3,
  output [31:0] io_out_bits_28_0,
  output [31:0] io_out_bits_28_1,
  output [31:0] io_out_bits_28_2,
  output [31:0] io_out_bits_28_3,
  output [31:0] io_out_bits_29_0,
  output [31:0] io_out_bits_29_1,
  output [31:0] io_out_bits_29_2,
  output [31:0] io_out_bits_29_3,
  output [31:0] io_out_bits_30_0,
  output [31:0] io_out_bits_30_1,
  output [31:0] io_out_bits_30_2,
  output [31:0] io_out_bits_30_3,
  output [31:0] io_out_bits_31_0,
  output [31:0] io_out_bits_31_1,
  output [31:0] io_out_bits_31_2,
  output [31:0] io_out_bits_31_3,
  output [31:0] io_out_bits_32_0,
  output [31:0] io_out_bits_32_1,
  output [31:0] io_out_bits_32_2,
  output [31:0] io_out_bits_32_3,
  output [31:0] io_out_bits_33_0,
  output [31:0] io_out_bits_33_1,
  output [31:0] io_out_bits_33_2,
  output [31:0] io_out_bits_33_3,
  output [31:0] io_out_bits_34_0,
  output [31:0] io_out_bits_34_1,
  output [31:0] io_out_bits_34_2,
  output [31:0] io_out_bits_34_3,
  output [31:0] io_out_bits_35_0,
  output [31:0] io_out_bits_35_1,
  output [31:0] io_out_bits_35_2,
  output [31:0] io_out_bits_35_3,
  output [31:0] io_out_bits_36_0,
  output [31:0] io_out_bits_36_1,
  output [31:0] io_out_bits_36_2,
  output [31:0] io_out_bits_36_3,
  output [31:0] io_out_bits_37_0,
  output [31:0] io_out_bits_37_1,
  output [31:0] io_out_bits_37_2,
  output [31:0] io_out_bits_37_3,
  output [31:0] io_out_bits_38_0,
  output [31:0] io_out_bits_38_1,
  output [31:0] io_out_bits_38_2,
  output [31:0] io_out_bits_38_3,
  output [31:0] io_out_bits_39_0,
  output [31:0] io_out_bits_39_1,
  output [31:0] io_out_bits_39_2,
  output [31:0] io_out_bits_39_3,
  output [31:0] io_out_bits_40_0,
  output [31:0] io_out_bits_40_1,
  output [31:0] io_out_bits_40_2,
  output [31:0] io_out_bits_40_3,
  output [31:0] io_out_bits_41_0,
  output [31:0] io_out_bits_41_1,
  output [31:0] io_out_bits_41_2,
  output [31:0] io_out_bits_41_3,
  output [31:0] io_out_bits_42_0,
  output [31:0] io_out_bits_42_1,
  output [31:0] io_out_bits_42_2,
  output [31:0] io_out_bits_42_3,
  output [31:0] io_out_bits_43_0,
  output [31:0] io_out_bits_43_1,
  output [31:0] io_out_bits_43_2,
  output [31:0] io_out_bits_43_3,
  output [31:0] io_out_bits_44_0,
  output [31:0] io_out_bits_44_1,
  output [31:0] io_out_bits_44_2,
  output [31:0] io_out_bits_44_3,
  output [31:0] io_out_bits_45_0,
  output [31:0] io_out_bits_45_1,
  output [31:0] io_out_bits_45_2,
  output [31:0] io_out_bits_45_3,
  output [31:0] io_out_bits_46_0,
  output [31:0] io_out_bits_46_1,
  output [31:0] io_out_bits_46_2,
  output [31:0] io_out_bits_46_3,
  output [31:0] io_out_bits_47_0,
  output [31:0] io_out_bits_47_1,
  output [31:0] io_out_bits_47_2,
  output [31:0] io_out_bits_47_3,
  output [31:0] io_out_bits_48_0,
  output [31:0] io_out_bits_48_1,
  output [31:0] io_out_bits_48_2,
  output [31:0] io_out_bits_48_3,
  output [31:0] io_out_bits_49_0,
  output [31:0] io_out_bits_49_1,
  output [31:0] io_out_bits_49_2,
  output [31:0] io_out_bits_49_3,
  output [31:0] io_out_bits_50_0,
  output [31:0] io_out_bits_50_1,
  output [31:0] io_out_bits_50_2,
  output [31:0] io_out_bits_50_3,
  output [31:0] io_out_bits_51_0,
  output [31:0] io_out_bits_51_1,
  output [31:0] io_out_bits_51_2,
  output [31:0] io_out_bits_51_3,
  output [31:0] io_out_bits_52_0,
  output [31:0] io_out_bits_52_1,
  output [31:0] io_out_bits_52_2,
  output [31:0] io_out_bits_52_3,
  output [31:0] io_out_bits_53_0,
  output [31:0] io_out_bits_53_1,
  output [31:0] io_out_bits_53_2,
  output [31:0] io_out_bits_53_3,
  output [31:0] io_out_bits_54_0,
  output [31:0] io_out_bits_54_1,
  output [31:0] io_out_bits_54_2,
  output [31:0] io_out_bits_54_3,
  output [31:0] io_out_bits_55_0,
  output [31:0] io_out_bits_55_1,
  output [31:0] io_out_bits_55_2,
  output [31:0] io_out_bits_55_3,
  output [31:0] io_out_bits_56_0,
  output [31:0] io_out_bits_56_1,
  output [31:0] io_out_bits_56_2,
  output [31:0] io_out_bits_56_3,
  output [31:0] io_out_bits_57_0,
  output [31:0] io_out_bits_57_1,
  output [31:0] io_out_bits_57_2,
  output [31:0] io_out_bits_57_3,
  output [31:0] io_out_bits_58_0,
  output [31:0] io_out_bits_58_1,
  output [31:0] io_out_bits_58_2,
  output [31:0] io_out_bits_58_3,
  output [31:0] io_out_bits_59_0,
  output [31:0] io_out_bits_59_1,
  output [31:0] io_out_bits_59_2,
  output [31:0] io_out_bits_59_3,
  output [31:0] io_out_bits_60_0,
  output [31:0] io_out_bits_60_1,
  output [31:0] io_out_bits_60_2,
  output [31:0] io_out_bits_60_3,
  output [31:0] io_out_bits_61_0,
  output [31:0] io_out_bits_61_1,
  output [31:0] io_out_bits_61_2,
  output [31:0] io_out_bits_61_3,
  output [31:0] io_out_bits_62_0,
  output [31:0] io_out_bits_62_1,
  output [31:0] io_out_bits_62_2,
  output [31:0] io_out_bits_62_3,
  output [31:0] io_out_bits_63_0,
  output [31:0] io_out_bits_63_1,
  output [31:0] io_out_bits_63_2,
  output [31:0] io_out_bits_63_3,
  output [31:0] io_out_bits_64_0,
  output [31:0] io_out_bits_64_1,
  output [31:0] io_out_bits_64_2,
  output [31:0] io_out_bits_64_3,
  output [31:0] io_out_bits_65_0,
  output [31:0] io_out_bits_65_1,
  output [31:0] io_out_bits_65_2,
  output [31:0] io_out_bits_65_3,
  output [31:0] io_out_bits_66_0,
  output [31:0] io_out_bits_66_1,
  output [31:0] io_out_bits_66_2,
  output [31:0] io_out_bits_66_3,
  output [31:0] io_out_bits_67_0,
  output [31:0] io_out_bits_67_1,
  output [31:0] io_out_bits_67_2,
  output [31:0] io_out_bits_67_3,
  output [31:0] io_out_bits_68_0,
  output [31:0] io_out_bits_68_1,
  output [31:0] io_out_bits_68_2,
  output [31:0] io_out_bits_68_3,
  output [31:0] io_out_bits_69_0,
  output [31:0] io_out_bits_69_1,
  output [31:0] io_out_bits_69_2,
  output [31:0] io_out_bits_69_3,
  output [31:0] io_out_bits_70_0,
  output [31:0] io_out_bits_70_1,
  output [31:0] io_out_bits_70_2,
  output [31:0] io_out_bits_70_3,
  output [31:0] io_out_bits_71_0,
  output [31:0] io_out_bits_71_1,
  output [31:0] io_out_bits_71_2,
  output [31:0] io_out_bits_71_3,
  output [31:0] io_out_bits_72_0,
  output [31:0] io_out_bits_72_1,
  output [31:0] io_out_bits_72_2,
  output [31:0] io_out_bits_72_3,
  output [31:0] io_out_bits_73_0,
  output [31:0] io_out_bits_73_1,
  output [31:0] io_out_bits_73_2,
  output [31:0] io_out_bits_73_3,
  output [31:0] io_out_bits_74_0,
  output [31:0] io_out_bits_74_1,
  output [31:0] io_out_bits_74_2,
  output [31:0] io_out_bits_74_3,
  output [31:0] io_out_bits_75_0,
  output [31:0] io_out_bits_75_1,
  output [31:0] io_out_bits_75_2,
  output [31:0] io_out_bits_75_3,
  output [31:0] io_out_bits_76_0,
  output [31:0] io_out_bits_76_1,
  output [31:0] io_out_bits_76_2,
  output [31:0] io_out_bits_76_3,
  output [31:0] io_out_bits_77_0,
  output [31:0] io_out_bits_77_1,
  output [31:0] io_out_bits_77_2,
  output [31:0] io_out_bits_77_3,
  output [31:0] io_out_bits_78_0,
  output [31:0] io_out_bits_78_1,
  output [31:0] io_out_bits_78_2,
  output [31:0] io_out_bits_78_3,
  output [31:0] io_out_bits_79_0,
  output [31:0] io_out_bits_79_1,
  output [31:0] io_out_bits_79_2,
  output [31:0] io_out_bits_79_3,
  output [31:0] io_out_bits_80_0,
  output [31:0] io_out_bits_80_1,
  output [31:0] io_out_bits_80_2,
  output [31:0] io_out_bits_80_3,
  output [31:0] io_out_bits_81_0,
  output [31:0] io_out_bits_81_1,
  output [31:0] io_out_bits_81_2,
  output [31:0] io_out_bits_81_3,
  output [31:0] io_out_bits_82_0,
  output [31:0] io_out_bits_82_1,
  output [31:0] io_out_bits_82_2,
  output [31:0] io_out_bits_82_3,
  output [31:0] io_out_bits_83_0,
  output [31:0] io_out_bits_83_1,
  output [31:0] io_out_bits_83_2,
  output [31:0] io_out_bits_83_3,
  output [31:0] io_out_bits_84_0,
  output [31:0] io_out_bits_84_1,
  output [31:0] io_out_bits_84_2,
  output [31:0] io_out_bits_84_3,
  output [31:0] io_out_bits_85_0,
  output [31:0] io_out_bits_85_1,
  output [31:0] io_out_bits_85_2,
  output [31:0] io_out_bits_85_3,
  output [31:0] io_out_bits_86_0,
  output [31:0] io_out_bits_86_1,
  output [31:0] io_out_bits_86_2,
  output [31:0] io_out_bits_86_3,
  output [31:0] io_out_bits_87_0,
  output [31:0] io_out_bits_87_1,
  output [31:0] io_out_bits_87_2,
  output [31:0] io_out_bits_87_3,
  output [31:0] io_out_bits_88_0,
  output [31:0] io_out_bits_88_1,
  output [31:0] io_out_bits_88_2,
  output [31:0] io_out_bits_88_3,
  output [31:0] io_out_bits_89_0,
  output [31:0] io_out_bits_89_1,
  output [31:0] io_out_bits_89_2,
  output [31:0] io_out_bits_89_3,
  output [31:0] io_out_bits_90_0,
  output [31:0] io_out_bits_90_1,
  output [31:0] io_out_bits_90_2,
  output [31:0] io_out_bits_90_3,
  output [31:0] io_out_bits_91_0,
  output [31:0] io_out_bits_91_1,
  output [31:0] io_out_bits_91_2,
  output [31:0] io_out_bits_91_3,
  output [31:0] io_out_bits_92_0,
  output [31:0] io_out_bits_92_1,
  output [31:0] io_out_bits_92_2,
  output [31:0] io_out_bits_92_3,
  output [31:0] io_out_bits_93_0,
  output [31:0] io_out_bits_93_1,
  output [31:0] io_out_bits_93_2,
  output [31:0] io_out_bits_93_3,
  output [31:0] io_out_bits_94_0,
  output [31:0] io_out_bits_94_1,
  output [31:0] io_out_bits_94_2,
  output [31:0] io_out_bits_94_3,
  output [31:0] io_out_bits_95_0,
  output [31:0] io_out_bits_95_1,
  output [31:0] io_out_bits_95_2,
  output [31:0] io_out_bits_95_3,
  output [31:0] io_out_bits_96_0,
  output [31:0] io_out_bits_96_1,
  output [31:0] io_out_bits_96_2,
  output [31:0] io_out_bits_96_3,
  output [31:0] io_out_bits_97_0,
  output [31:0] io_out_bits_97_1,
  output [31:0] io_out_bits_97_2,
  output [31:0] io_out_bits_97_3,
  output [31:0] io_out_bits_98_0,
  output [31:0] io_out_bits_98_1,
  output [31:0] io_out_bits_98_2,
  output [31:0] io_out_bits_98_3,
  output [31:0] io_out_bits_99_0,
  output [31:0] io_out_bits_99_1,
  output [31:0] io_out_bits_99_2,
  output [31:0] io_out_bits_99_3
);
  reg [31:0] regs_0; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_0;
  reg [31:0] regs_1; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_1;
  reg [31:0] regs_2; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_2;
  reg [31:0] regs_3; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_3;
  reg [31:0] regs_4; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_4;
  reg [31:0] regs_5; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_5;
  reg [31:0] regs_6; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_6;
  reg [31:0] regs_7; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_7;
  reg [31:0] regs_8; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_8;
  reg [31:0] regs_9; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_9;
  reg [31:0] regs_10; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_10;
  reg [31:0] regs_11; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_11;
  reg [31:0] regs_12; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_12;
  reg [31:0] regs_13; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_13;
  reg [31:0] regs_14; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_14;
  reg [31:0] regs_15; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_15;
  reg [31:0] regs_16; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_16;
  reg [31:0] regs_17; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_17;
  reg [31:0] regs_18; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_18;
  reg [31:0] regs_19; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_19;
  reg [31:0] regs_20; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_20;
  reg [31:0] regs_21; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_21;
  reg [31:0] regs_22; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_22;
  reg [31:0] regs_23; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_23;
  reg [31:0] regs_24; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_24;
  reg [31:0] regs_25; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_25;
  reg [31:0] regs_26; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_26;
  reg [31:0] regs_27; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_27;
  reg [31:0] regs_28; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_28;
  reg [31:0] regs_29; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_29;
  reg [31:0] regs_30; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_30;
  reg [31:0] regs_31; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_31;
  reg [31:0] regs_32; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_32;
  reg [31:0] regs_33; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_33;
  reg [31:0] regs_34; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_34;
  reg [31:0] regs_35; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_35;
  reg [31:0] regs_36; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_36;
  reg [31:0] regs_37; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_37;
  reg [31:0] regs_38; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_38;
  reg [31:0] regs_39; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_39;
  reg [31:0] regs_40; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_40;
  reg [31:0] regs_41; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_41;
  reg [31:0] regs_42; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_42;
  reg [31:0] regs_43; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_43;
  reg [31:0] regs_44; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_44;
  reg [31:0] regs_45; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_45;
  reg [31:0] regs_46; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_46;
  reg [31:0] regs_47; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_47;
  reg [31:0] regs_48; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_48;
  reg [31:0] regs_49; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_49;
  reg [31:0] regs_50; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_50;
  reg [31:0] regs_51; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_51;
  reg [31:0] regs_52; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_52;
  reg [31:0] regs_53; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_53;
  reg [31:0] regs_54; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_54;
  reg [31:0] regs_55; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_55;
  reg [31:0] regs_56; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_56;
  reg [31:0] regs_57; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_57;
  reg [31:0] regs_58; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_58;
  reg [31:0] regs_59; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_59;
  reg [31:0] regs_60; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_60;
  reg [31:0] regs_61; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_61;
  reg [31:0] regs_62; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_62;
  reg [31:0] regs_63; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_63;
  reg [31:0] regs_64; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_64;
  reg [31:0] regs_65; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_65;
  reg [31:0] regs_66; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_66;
  reg [31:0] regs_67; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_67;
  reg [31:0] regs_68; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_68;
  reg [31:0] regs_69; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_69;
  reg [31:0] regs_70; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_70;
  reg [31:0] regs_71; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_71;
  reg [31:0] regs_72; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_72;
  reg [31:0] regs_73; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_73;
  reg [31:0] regs_74; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_74;
  reg [31:0] regs_75; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_75;
  reg [31:0] regs_76; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_76;
  reg [31:0] regs_77; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_77;
  reg [31:0] regs_78; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_78;
  reg [31:0] regs_79; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_79;
  reg [31:0] regs_80; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_80;
  reg [31:0] regs_81; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_81;
  reg [31:0] regs_82; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_82;
  reg [31:0] regs_83; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_83;
  reg [31:0] regs_84; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_84;
  reg [31:0] regs_85; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_85;
  reg [31:0] regs_86; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_86;
  reg [31:0] regs_87; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_87;
  reg [31:0] regs_88; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_88;
  reg [31:0] regs_89; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_89;
  reg [31:0] regs_90; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_90;
  reg [31:0] regs_91; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_91;
  reg [31:0] regs_92; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_92;
  reg [31:0] regs_93; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_93;
  reg [31:0] regs_94; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_94;
  reg [31:0] regs_95; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_95;
  reg [31:0] regs_96; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_96;
  reg [31:0] regs_97; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_97;
  reg [31:0] regs_98; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_98;
  reg [31:0] regs_99; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_99;
  reg [31:0] regs_100; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_100;
  reg [31:0] regs_101; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_101;
  reg [31:0] regs_102; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_102;
  reg [31:0] regs_103; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_103;
  reg [31:0] regs_104; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_104;
  reg [31:0] regs_105; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_105;
  reg [31:0] regs_106; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_106;
  reg [31:0] regs_107; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_107;
  reg [31:0] regs_108; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_108;
  reg [31:0] regs_109; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_109;
  reg [31:0] regs_110; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_110;
  reg [31:0] regs_111; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_111;
  reg [31:0] regs_112; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_112;
  reg [31:0] regs_113; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_113;
  reg [31:0] regs_114; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_114;
  reg [31:0] regs_115; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_115;
  reg [31:0] regs_116; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_116;
  reg [31:0] regs_117; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_117;
  reg [31:0] regs_118; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_118;
  reg [31:0] regs_119; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_119;
  reg [31:0] regs_120; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_120;
  reg [31:0] regs_121; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_121;
  reg [31:0] regs_122; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_122;
  reg [31:0] regs_123; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_123;
  reg [31:0] regs_124; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_124;
  reg [31:0] regs_125; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_125;
  reg [31:0] regs_126; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_126;
  reg [31:0] regs_127; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_127;
  reg [31:0] regs_128; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_128;
  reg [31:0] regs_129; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_129;
  reg [31:0] regs_130; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_130;
  reg [31:0] regs_131; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_131;
  reg [31:0] regs_132; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_132;
  reg [31:0] regs_133; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_133;
  reg [31:0] regs_134; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_134;
  reg [31:0] regs_135; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_135;
  reg [31:0] regs_136; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_136;
  reg [31:0] regs_137; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_137;
  reg [31:0] regs_138; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_138;
  reg [31:0] regs_139; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_139;
  reg [31:0] regs_140; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_140;
  reg [31:0] regs_141; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_141;
  reg [31:0] regs_142; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_142;
  reg [31:0] regs_143; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_143;
  reg [31:0] regs_144; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_144;
  reg [31:0] regs_145; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_145;
  reg [31:0] regs_146; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_146;
  reg [31:0] regs_147; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_147;
  reg [31:0] regs_148; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_148;
  reg [31:0] regs_149; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_149;
  reg [31:0] regs_150; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_150;
  reg [31:0] regs_151; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_151;
  reg [31:0] regs_152; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_152;
  reg [31:0] regs_153; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_153;
  reg [31:0] regs_154; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_154;
  reg [31:0] regs_155; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_155;
  reg [31:0] regs_156; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_156;
  reg [31:0] regs_157; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_157;
  reg [31:0] regs_158; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_158;
  reg [31:0] regs_159; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_159;
  reg [31:0] regs_160; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_160;
  reg [31:0] regs_161; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_161;
  reg [31:0] regs_162; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_162;
  reg [31:0] regs_163; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_163;
  reg [31:0] regs_164; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_164;
  reg [31:0] regs_165; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_165;
  reg [31:0] regs_166; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_166;
  reg [31:0] regs_167; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_167;
  reg [31:0] regs_168; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_168;
  reg [31:0] regs_169; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_169;
  reg [31:0] regs_170; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_170;
  reg [31:0] regs_171; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_171;
  reg [31:0] regs_172; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_172;
  reg [31:0] regs_173; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_173;
  reg [31:0] regs_174; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_174;
  reg [31:0] regs_175; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_175;
  reg [31:0] regs_176; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_176;
  reg [31:0] regs_177; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_177;
  reg [31:0] regs_178; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_178;
  reg [31:0] regs_179; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_179;
  reg [31:0] regs_180; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_180;
  reg [31:0] regs_181; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_181;
  reg [31:0] regs_182; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_182;
  reg [31:0] regs_183; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_183;
  reg [31:0] regs_184; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_184;
  reg [31:0] regs_185; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_185;
  reg [31:0] regs_186; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_186;
  reg [31:0] regs_187; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_187;
  reg [31:0] regs_188; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_188;
  reg [31:0] regs_189; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_189;
  reg [31:0] regs_190; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_190;
  reg [31:0] regs_191; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_191;
  reg [31:0] regs_192; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_192;
  reg [31:0] regs_193; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_193;
  reg [31:0] regs_194; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_194;
  reg [31:0] regs_195; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_195;
  reg [31:0] regs_196; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_196;
  reg [31:0] regs_197; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_197;
  reg [31:0] regs_198; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_198;
  reg [31:0] regs_199; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_199;
  reg [31:0] regs_200; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_200;
  reg [31:0] regs_201; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_201;
  reg [31:0] regs_202; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_202;
  reg [31:0] regs_203; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_203;
  reg [31:0] regs_204; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_204;
  reg [31:0] regs_205; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_205;
  reg [31:0] regs_206; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_206;
  reg [31:0] regs_207; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_207;
  reg [31:0] regs_208; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_208;
  reg [31:0] regs_209; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_209;
  reg [31:0] regs_210; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_210;
  reg [31:0] regs_211; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_211;
  reg [31:0] regs_212; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_212;
  reg [31:0] regs_213; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_213;
  reg [31:0] regs_214; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_214;
  reg [31:0] regs_215; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_215;
  reg [31:0] regs_216; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_216;
  reg [31:0] regs_217; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_217;
  reg [31:0] regs_218; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_218;
  reg [31:0] regs_219; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_219;
  reg [31:0] regs_220; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_220;
  reg [31:0] regs_221; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_221;
  reg [31:0] regs_222; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_222;
  reg [31:0] regs_223; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_223;
  reg [31:0] regs_224; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_224;
  reg [31:0] regs_225; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_225;
  reg [31:0] regs_226; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_226;
  reg [31:0] regs_227; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_227;
  reg [31:0] regs_228; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_228;
  reg [31:0] regs_229; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_229;
  reg [31:0] regs_230; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_230;
  reg [31:0] regs_231; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_231;
  reg [31:0] regs_232; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_232;
  reg [31:0] regs_233; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_233;
  reg [31:0] regs_234; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_234;
  reg [31:0] regs_235; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_235;
  reg [31:0] regs_236; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_236;
  reg [31:0] regs_237; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_237;
  reg [31:0] regs_238; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_238;
  reg [31:0] regs_239; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_239;
  reg [31:0] regs_240; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_240;
  reg [31:0] regs_241; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_241;
  reg [31:0] regs_242; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_242;
  reg [31:0] regs_243; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_243;
  reg [31:0] regs_244; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_244;
  reg [31:0] regs_245; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_245;
  reg [31:0] regs_246; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_246;
  reg [31:0] regs_247; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_247;
  reg [31:0] regs_248; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_248;
  reg [31:0] regs_249; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_249;
  reg [31:0] regs_250; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_250;
  reg [31:0] regs_251; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_251;
  reg [31:0] regs_252; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_252;
  reg [31:0] regs_253; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_253;
  reg [31:0] regs_254; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_254;
  reg [31:0] regs_255; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_255;
  reg [31:0] regs_256; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_256;
  reg [31:0] regs_257; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_257;
  reg [31:0] regs_258; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_258;
  reg [31:0] regs_259; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_259;
  reg [31:0] regs_260; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_260;
  reg [31:0] regs_261; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_261;
  reg [31:0] regs_262; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_262;
  reg [31:0] regs_263; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_263;
  reg [31:0] regs_264; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_264;
  reg [31:0] regs_265; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_265;
  reg [31:0] regs_266; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_266;
  reg [31:0] regs_267; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_267;
  reg [31:0] regs_268; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_268;
  reg [31:0] regs_269; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_269;
  reg [31:0] regs_270; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_270;
  reg [31:0] regs_271; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_271;
  reg [31:0] regs_272; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_272;
  reg [31:0] regs_273; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_273;
  reg [31:0] regs_274; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_274;
  reg [31:0] regs_275; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_275;
  reg [31:0] regs_276; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_276;
  reg [31:0] regs_277; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_277;
  reg [31:0] regs_278; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_278;
  reg [31:0] regs_279; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_279;
  reg [31:0] regs_280; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_280;
  reg [31:0] regs_281; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_281;
  reg [31:0] regs_282; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_282;
  reg [31:0] regs_283; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_283;
  reg [31:0] regs_284; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_284;
  reg [31:0] regs_285; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_285;
  reg [31:0] regs_286; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_286;
  reg [31:0] regs_287; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_287;
  reg [31:0] regs_288; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_288;
  reg [31:0] regs_289; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_289;
  reg [31:0] regs_290; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_290;
  reg [31:0] regs_291; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_291;
  reg [31:0] regs_292; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_292;
  reg [31:0] regs_293; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_293;
  reg [31:0] regs_294; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_294;
  reg [31:0] regs_295; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_295;
  reg [31:0] regs_296; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_296;
  reg [31:0] regs_297; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_297;
  reg [31:0] regs_298; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_298;
  reg [31:0] regs_299; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_299;
  reg [31:0] regs_300; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_300;
  reg [31:0] regs_301; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_301;
  reg [31:0] regs_302; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_302;
  reg [31:0] regs_303; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_303;
  reg [31:0] regs_304; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_304;
  reg [31:0] regs_305; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_305;
  reg [31:0] regs_306; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_306;
  reg [31:0] regs_307; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_307;
  reg [31:0] regs_308; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_308;
  reg [31:0] regs_309; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_309;
  reg [31:0] regs_310; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_310;
  reg [31:0] regs_311; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_311;
  reg [31:0] regs_312; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_312;
  reg [31:0] regs_313; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_313;
  reg [31:0] regs_314; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_314;
  reg [31:0] regs_315; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_315;
  reg [31:0] regs_316; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_316;
  reg [31:0] regs_317; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_317;
  reg [31:0] regs_318; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_318;
  reg [31:0] regs_319; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_319;
  reg [31:0] regs_320; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_320;
  reg [31:0] regs_321; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_321;
  reg [31:0] regs_322; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_322;
  reg [31:0] regs_323; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_323;
  reg [31:0] regs_324; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_324;
  reg [31:0] regs_325; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_325;
  reg [31:0] regs_326; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_326;
  reg [31:0] regs_327; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_327;
  reg [31:0] regs_328; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_328;
  reg [31:0] regs_329; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_329;
  reg [31:0] regs_330; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_330;
  reg [31:0] regs_331; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_331;
  reg [31:0] regs_332; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_332;
  reg [31:0] regs_333; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_333;
  reg [31:0] regs_334; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_334;
  reg [31:0] regs_335; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_335;
  reg [31:0] regs_336; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_336;
  reg [31:0] regs_337; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_337;
  reg [31:0] regs_338; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_338;
  reg [31:0] regs_339; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_339;
  reg [31:0] regs_340; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_340;
  reg [31:0] regs_341; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_341;
  reg [31:0] regs_342; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_342;
  reg [31:0] regs_343; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_343;
  reg [31:0] regs_344; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_344;
  reg [31:0] regs_345; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_345;
  reg [31:0] regs_346; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_346;
  reg [31:0] regs_347; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_347;
  reg [31:0] regs_348; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_348;
  reg [31:0] regs_349; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_349;
  reg [31:0] regs_350; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_350;
  reg [31:0] regs_351; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_351;
  reg [31:0] regs_352; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_352;
  reg [31:0] regs_353; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_353;
  reg [31:0] regs_354; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_354;
  reg [31:0] regs_355; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_355;
  reg [31:0] regs_356; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_356;
  reg [31:0] regs_357; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_357;
  reg [31:0] regs_358; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_358;
  reg [31:0] regs_359; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_359;
  reg [31:0] regs_360; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_360;
  reg [31:0] regs_361; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_361;
  reg [31:0] regs_362; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_362;
  reg [31:0] regs_363; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_363;
  reg [31:0] regs_364; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_364;
  reg [31:0] regs_365; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_365;
  reg [31:0] regs_366; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_366;
  reg [31:0] regs_367; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_367;
  reg [31:0] regs_368; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_368;
  reg [31:0] regs_369; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_369;
  reg [31:0] regs_370; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_370;
  reg [31:0] regs_371; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_371;
  reg [31:0] regs_372; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_372;
  reg [31:0] regs_373; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_373;
  reg [31:0] regs_374; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_374;
  reg [31:0] regs_375; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_375;
  reg [31:0] regs_376; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_376;
  reg [31:0] regs_377; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_377;
  reg [31:0] regs_378; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_378;
  reg [31:0] regs_379; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_379;
  reg [31:0] regs_380; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_380;
  reg [31:0] regs_381; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_381;
  reg [31:0] regs_382; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_382;
  reg [31:0] regs_383; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_383;
  reg [31:0] regs_384; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_384;
  reg [31:0] regs_385; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_385;
  reg [31:0] regs_386; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_386;
  reg [31:0] regs_387; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_387;
  reg [31:0] regs_388; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_388;
  reg [31:0] regs_389; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_389;
  reg [31:0] regs_390; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_390;
  reg [31:0] regs_391; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_391;
  reg [31:0] regs_392; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_392;
  reg [31:0] regs_393; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_393;
  reg [31:0] regs_394; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_394;
  reg [31:0] regs_395; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_395;
  reg [31:0] regs_396; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_396;
  reg [31:0] regs_397; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_397;
  reg [31:0] regs_398; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_398;
  reg [31:0] regs_399; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_399;
  assign io_out_bits_0_0 = regs_0; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_1 = regs_1; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_2 = regs_2; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_3 = regs_3; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_1_0 = regs_4; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_1_1 = regs_5; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_1_2 = regs_6; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_1_3 = regs_7; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_2_0 = regs_8; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_2_1 = regs_9; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_2_2 = regs_10; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_2_3 = regs_11; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_3_0 = regs_12; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_3_1 = regs_13; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_3_2 = regs_14; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_3_3 = regs_15; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_4_0 = regs_16; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_4_1 = regs_17; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_4_2 = regs_18; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_4_3 = regs_19; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_5_0 = regs_20; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_5_1 = regs_21; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_5_2 = regs_22; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_5_3 = regs_23; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_6_0 = regs_24; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_6_1 = regs_25; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_6_2 = regs_26; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_6_3 = regs_27; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_7_0 = regs_28; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_7_1 = regs_29; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_7_2 = regs_30; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_7_3 = regs_31; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_8_0 = regs_32; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_8_1 = regs_33; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_8_2 = regs_34; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_8_3 = regs_35; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_9_0 = regs_36; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_9_1 = regs_37; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_9_2 = regs_38; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_9_3 = regs_39; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_10_0 = regs_40; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_10_1 = regs_41; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_10_2 = regs_42; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_10_3 = regs_43; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_11_0 = regs_44; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_11_1 = regs_45; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_11_2 = regs_46; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_11_3 = regs_47; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_12_0 = regs_48; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_12_1 = regs_49; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_12_2 = regs_50; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_12_3 = regs_51; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_13_0 = regs_52; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_13_1 = regs_53; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_13_2 = regs_54; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_13_3 = regs_55; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_14_0 = regs_56; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_14_1 = regs_57; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_14_2 = regs_58; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_14_3 = regs_59; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_15_0 = regs_60; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_15_1 = regs_61; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_15_2 = regs_62; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_15_3 = regs_63; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_16_0 = regs_64; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_16_1 = regs_65; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_16_2 = regs_66; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_16_3 = regs_67; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_17_0 = regs_68; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_17_1 = regs_69; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_17_2 = regs_70; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_17_3 = regs_71; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_18_0 = regs_72; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_18_1 = regs_73; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_18_2 = regs_74; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_18_3 = regs_75; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_19_0 = regs_76; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_19_1 = regs_77; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_19_2 = regs_78; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_19_3 = regs_79; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_20_0 = regs_80; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_20_1 = regs_81; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_20_2 = regs_82; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_20_3 = regs_83; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_21_0 = regs_84; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_21_1 = regs_85; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_21_2 = regs_86; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_21_3 = regs_87; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_22_0 = regs_88; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_22_1 = regs_89; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_22_2 = regs_90; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_22_3 = regs_91; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_23_0 = regs_92; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_23_1 = regs_93; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_23_2 = regs_94; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_23_3 = regs_95; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_24_0 = regs_96; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_24_1 = regs_97; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_24_2 = regs_98; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_24_3 = regs_99; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_25_0 = regs_100; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_25_1 = regs_101; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_25_2 = regs_102; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_25_3 = regs_103; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_26_0 = regs_104; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_26_1 = regs_105; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_26_2 = regs_106; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_26_3 = regs_107; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_27_0 = regs_108; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_27_1 = regs_109; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_27_2 = regs_110; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_27_3 = regs_111; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_28_0 = regs_112; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_28_1 = regs_113; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_28_2 = regs_114; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_28_3 = regs_115; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_29_0 = regs_116; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_29_1 = regs_117; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_29_2 = regs_118; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_29_3 = regs_119; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_30_0 = regs_120; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_30_1 = regs_121; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_30_2 = regs_122; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_30_3 = regs_123; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_31_0 = regs_124; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_31_1 = regs_125; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_31_2 = regs_126; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_31_3 = regs_127; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_32_0 = regs_128; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_32_1 = regs_129; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_32_2 = regs_130; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_32_3 = regs_131; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_33_0 = regs_132; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_33_1 = regs_133; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_33_2 = regs_134; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_33_3 = regs_135; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_34_0 = regs_136; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_34_1 = regs_137; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_34_2 = regs_138; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_34_3 = regs_139; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_35_0 = regs_140; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_35_1 = regs_141; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_35_2 = regs_142; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_35_3 = regs_143; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_36_0 = regs_144; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_36_1 = regs_145; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_36_2 = regs_146; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_36_3 = regs_147; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_37_0 = regs_148; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_37_1 = regs_149; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_37_2 = regs_150; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_37_3 = regs_151; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_38_0 = regs_152; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_38_1 = regs_153; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_38_2 = regs_154; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_38_3 = regs_155; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_39_0 = regs_156; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_39_1 = regs_157; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_39_2 = regs_158; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_39_3 = regs_159; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_40_0 = regs_160; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_40_1 = regs_161; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_40_2 = regs_162; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_40_3 = regs_163; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_41_0 = regs_164; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_41_1 = regs_165; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_41_2 = regs_166; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_41_3 = regs_167; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_42_0 = regs_168; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_42_1 = regs_169; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_42_2 = regs_170; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_42_3 = regs_171; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_43_0 = regs_172; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_43_1 = regs_173; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_43_2 = regs_174; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_43_3 = regs_175; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_44_0 = regs_176; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_44_1 = regs_177; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_44_2 = regs_178; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_44_3 = regs_179; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_45_0 = regs_180; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_45_1 = regs_181; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_45_2 = regs_182; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_45_3 = regs_183; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_46_0 = regs_184; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_46_1 = regs_185; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_46_2 = regs_186; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_46_3 = regs_187; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_47_0 = regs_188; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_47_1 = regs_189; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_47_2 = regs_190; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_47_3 = regs_191; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_48_0 = regs_192; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_48_1 = regs_193; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_48_2 = regs_194; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_48_3 = regs_195; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_49_0 = regs_196; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_49_1 = regs_197; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_49_2 = regs_198; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_49_3 = regs_199; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_50_0 = regs_200; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_50_1 = regs_201; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_50_2 = regs_202; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_50_3 = regs_203; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_51_0 = regs_204; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_51_1 = regs_205; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_51_2 = regs_206; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_51_3 = regs_207; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_52_0 = regs_208; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_52_1 = regs_209; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_52_2 = regs_210; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_52_3 = regs_211; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_53_0 = regs_212; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_53_1 = regs_213; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_53_2 = regs_214; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_53_3 = regs_215; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_54_0 = regs_216; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_54_1 = regs_217; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_54_2 = regs_218; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_54_3 = regs_219; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_55_0 = regs_220; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_55_1 = regs_221; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_55_2 = regs_222; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_55_3 = regs_223; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_56_0 = regs_224; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_56_1 = regs_225; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_56_2 = regs_226; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_56_3 = regs_227; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_57_0 = regs_228; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_57_1 = regs_229; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_57_2 = regs_230; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_57_3 = regs_231; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_58_0 = regs_232; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_58_1 = regs_233; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_58_2 = regs_234; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_58_3 = regs_235; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_59_0 = regs_236; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_59_1 = regs_237; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_59_2 = regs_238; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_59_3 = regs_239; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_60_0 = regs_240; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_60_1 = regs_241; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_60_2 = regs_242; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_60_3 = regs_243; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_61_0 = regs_244; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_61_1 = regs_245; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_61_2 = regs_246; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_61_3 = regs_247; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_62_0 = regs_248; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_62_1 = regs_249; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_62_2 = regs_250; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_62_3 = regs_251; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_63_0 = regs_252; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_63_1 = regs_253; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_63_2 = regs_254; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_63_3 = regs_255; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_64_0 = regs_256; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_64_1 = regs_257; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_64_2 = regs_258; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_64_3 = regs_259; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_65_0 = regs_260; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_65_1 = regs_261; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_65_2 = regs_262; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_65_3 = regs_263; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_66_0 = regs_264; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_66_1 = regs_265; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_66_2 = regs_266; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_66_3 = regs_267; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_67_0 = regs_268; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_67_1 = regs_269; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_67_2 = regs_270; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_67_3 = regs_271; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_68_0 = regs_272; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_68_1 = regs_273; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_68_2 = regs_274; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_68_3 = regs_275; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_69_0 = regs_276; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_69_1 = regs_277; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_69_2 = regs_278; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_69_3 = regs_279; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_70_0 = regs_280; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_70_1 = regs_281; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_70_2 = regs_282; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_70_3 = regs_283; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_71_0 = regs_284; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_71_1 = regs_285; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_71_2 = regs_286; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_71_3 = regs_287; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_72_0 = regs_288; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_72_1 = regs_289; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_72_2 = regs_290; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_72_3 = regs_291; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_73_0 = regs_292; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_73_1 = regs_293; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_73_2 = regs_294; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_73_3 = regs_295; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_74_0 = regs_296; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_74_1 = regs_297; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_74_2 = regs_298; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_74_3 = regs_299; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_75_0 = regs_300; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_75_1 = regs_301; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_75_2 = regs_302; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_75_3 = regs_303; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_76_0 = regs_304; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_76_1 = regs_305; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_76_2 = regs_306; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_76_3 = regs_307; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_77_0 = regs_308; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_77_1 = regs_309; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_77_2 = regs_310; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_77_3 = regs_311; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_78_0 = regs_312; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_78_1 = regs_313; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_78_2 = regs_314; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_78_3 = regs_315; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_79_0 = regs_316; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_79_1 = regs_317; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_79_2 = regs_318; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_79_3 = regs_319; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_80_0 = regs_320; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_80_1 = regs_321; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_80_2 = regs_322; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_80_3 = regs_323; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_81_0 = regs_324; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_81_1 = regs_325; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_81_2 = regs_326; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_81_3 = regs_327; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_82_0 = regs_328; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_82_1 = regs_329; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_82_2 = regs_330; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_82_3 = regs_331; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_83_0 = regs_332; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_83_1 = regs_333; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_83_2 = regs_334; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_83_3 = regs_335; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_84_0 = regs_336; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_84_1 = regs_337; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_84_2 = regs_338; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_84_3 = regs_339; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_85_0 = regs_340; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_85_1 = regs_341; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_85_2 = regs_342; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_85_3 = regs_343; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_86_0 = regs_344; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_86_1 = regs_345; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_86_2 = regs_346; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_86_3 = regs_347; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_87_0 = regs_348; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_87_1 = regs_349; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_87_2 = regs_350; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_87_3 = regs_351; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_88_0 = regs_352; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_88_1 = regs_353; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_88_2 = regs_354; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_88_3 = regs_355; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_89_0 = regs_356; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_89_1 = regs_357; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_89_2 = regs_358; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_89_3 = regs_359; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_90_0 = regs_360; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_90_1 = regs_361; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_90_2 = regs_362; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_90_3 = regs_363; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_91_0 = regs_364; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_91_1 = regs_365; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_91_2 = regs_366; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_91_3 = regs_367; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_92_0 = regs_368; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_92_1 = regs_369; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_92_2 = regs_370; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_92_3 = regs_371; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_93_0 = regs_372; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_93_1 = regs_373; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_93_2 = regs_374; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_93_3 = regs_375; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_94_0 = regs_376; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_94_1 = regs_377; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_94_2 = regs_378; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_94_3 = regs_379; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_95_0 = regs_380; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_95_1 = regs_381; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_95_2 = regs_382; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_95_3 = regs_383; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_96_0 = regs_384; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_96_1 = regs_385; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_96_2 = regs_386; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_96_3 = regs_387; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_97_0 = regs_388; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_97_1 = regs_389; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_97_2 = regs_390; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_97_3 = regs_391; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_98_0 = regs_392; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_98_1 = regs_393; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_98_2 = regs_394; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_98_3 = regs_395; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_99_0 = regs_396; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_99_1 = regs_397; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_99_2 = regs_398; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_99_3 = regs_399; // @[MemoryBuffer.scala 65:25]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  regs_3 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  regs_4 = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  regs_5 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  regs_6 = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  regs_7 = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  regs_8 = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  regs_9 = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  regs_10 = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  regs_11 = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  regs_12 = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  regs_13 = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  regs_14 = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  regs_15 = _RAND_15[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  regs_16 = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  regs_17 = _RAND_17[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  regs_18 = _RAND_18[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  regs_19 = _RAND_19[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  regs_20 = _RAND_20[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  regs_21 = _RAND_21[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  regs_22 = _RAND_22[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  regs_23 = _RAND_23[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  regs_24 = _RAND_24[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  regs_25 = _RAND_25[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  regs_26 = _RAND_26[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  regs_27 = _RAND_27[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  regs_28 = _RAND_28[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  regs_29 = _RAND_29[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  regs_30 = _RAND_30[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  regs_31 = _RAND_31[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  regs_32 = _RAND_32[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  regs_33 = _RAND_33[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  regs_34 = _RAND_34[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  regs_35 = _RAND_35[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  regs_36 = _RAND_36[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  regs_37 = _RAND_37[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  regs_38 = _RAND_38[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  regs_39 = _RAND_39[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  regs_40 = _RAND_40[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  regs_41 = _RAND_41[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  regs_42 = _RAND_42[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  regs_43 = _RAND_43[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  regs_44 = _RAND_44[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  regs_45 = _RAND_45[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  regs_46 = _RAND_46[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  regs_47 = _RAND_47[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  regs_48 = _RAND_48[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  regs_49 = _RAND_49[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  regs_50 = _RAND_50[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  regs_51 = _RAND_51[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  regs_52 = _RAND_52[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  regs_53 = _RAND_53[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  regs_54 = _RAND_54[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  regs_55 = _RAND_55[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  regs_56 = _RAND_56[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  regs_57 = _RAND_57[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  regs_58 = _RAND_58[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  regs_59 = _RAND_59[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  regs_60 = _RAND_60[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  regs_61 = _RAND_61[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  regs_62 = _RAND_62[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  regs_63 = _RAND_63[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  regs_64 = _RAND_64[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  regs_65 = _RAND_65[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  regs_66 = _RAND_66[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  regs_67 = _RAND_67[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  regs_68 = _RAND_68[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  regs_69 = _RAND_69[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  regs_70 = _RAND_70[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  regs_71 = _RAND_71[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  regs_72 = _RAND_72[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  regs_73 = _RAND_73[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  regs_74 = _RAND_74[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  regs_75 = _RAND_75[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  regs_76 = _RAND_76[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  regs_77 = _RAND_77[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  regs_78 = _RAND_78[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  regs_79 = _RAND_79[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  regs_80 = _RAND_80[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  regs_81 = _RAND_81[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  regs_82 = _RAND_82[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  regs_83 = _RAND_83[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  regs_84 = _RAND_84[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  regs_85 = _RAND_85[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  regs_86 = _RAND_86[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  regs_87 = _RAND_87[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  regs_88 = _RAND_88[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  regs_89 = _RAND_89[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  regs_90 = _RAND_90[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  regs_91 = _RAND_91[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  regs_92 = _RAND_92[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  regs_93 = _RAND_93[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  regs_94 = _RAND_94[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  regs_95 = _RAND_95[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  regs_96 = _RAND_96[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  regs_97 = _RAND_97[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  regs_98 = _RAND_98[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  regs_99 = _RAND_99[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  regs_100 = _RAND_100[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  regs_101 = _RAND_101[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  regs_102 = _RAND_102[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  regs_103 = _RAND_103[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  regs_104 = _RAND_104[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  regs_105 = _RAND_105[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  regs_106 = _RAND_106[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  regs_107 = _RAND_107[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  regs_108 = _RAND_108[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  regs_109 = _RAND_109[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  regs_110 = _RAND_110[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  regs_111 = _RAND_111[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  regs_112 = _RAND_112[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  regs_113 = _RAND_113[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  regs_114 = _RAND_114[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  regs_115 = _RAND_115[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  regs_116 = _RAND_116[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  regs_117 = _RAND_117[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  regs_118 = _RAND_118[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  regs_119 = _RAND_119[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  regs_120 = _RAND_120[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  regs_121 = _RAND_121[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  regs_122 = _RAND_122[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  regs_123 = _RAND_123[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  regs_124 = _RAND_124[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  regs_125 = _RAND_125[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  regs_126 = _RAND_126[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  regs_127 = _RAND_127[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  regs_128 = _RAND_128[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  regs_129 = _RAND_129[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  regs_130 = _RAND_130[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  regs_131 = _RAND_131[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  regs_132 = _RAND_132[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  regs_133 = _RAND_133[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  regs_134 = _RAND_134[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  regs_135 = _RAND_135[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  regs_136 = _RAND_136[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  regs_137 = _RAND_137[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  regs_138 = _RAND_138[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  regs_139 = _RAND_139[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  regs_140 = _RAND_140[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  regs_141 = _RAND_141[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  regs_142 = _RAND_142[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  regs_143 = _RAND_143[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  regs_144 = _RAND_144[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  regs_145 = _RAND_145[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  regs_146 = _RAND_146[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{`RANDOM}};
  regs_147 = _RAND_147[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{`RANDOM}};
  regs_148 = _RAND_148[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{`RANDOM}};
  regs_149 = _RAND_149[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{`RANDOM}};
  regs_150 = _RAND_150[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{`RANDOM}};
  regs_151 = _RAND_151[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{`RANDOM}};
  regs_152 = _RAND_152[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  regs_153 = _RAND_153[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  regs_154 = _RAND_154[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  regs_155 = _RAND_155[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  regs_156 = _RAND_156[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  regs_157 = _RAND_157[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  regs_158 = _RAND_158[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  regs_159 = _RAND_159[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  regs_160 = _RAND_160[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  regs_161 = _RAND_161[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  regs_162 = _RAND_162[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  regs_163 = _RAND_163[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  regs_164 = _RAND_164[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  regs_165 = _RAND_165[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  regs_166 = _RAND_166[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  regs_167 = _RAND_167[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  regs_168 = _RAND_168[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{`RANDOM}};
  regs_169 = _RAND_169[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{`RANDOM}};
  regs_170 = _RAND_170[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  regs_171 = _RAND_171[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  regs_172 = _RAND_172[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{`RANDOM}};
  regs_173 = _RAND_173[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  regs_174 = _RAND_174[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  regs_175 = _RAND_175[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  regs_176 = _RAND_176[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  regs_177 = _RAND_177[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  regs_178 = _RAND_178[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{`RANDOM}};
  regs_179 = _RAND_179[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  regs_180 = _RAND_180[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{`RANDOM}};
  regs_181 = _RAND_181[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  regs_182 = _RAND_182[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  regs_183 = _RAND_183[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  regs_184 = _RAND_184[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  regs_185 = _RAND_185[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  regs_186 = _RAND_186[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  regs_187 = _RAND_187[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  regs_188 = _RAND_188[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{`RANDOM}};
  regs_189 = _RAND_189[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{`RANDOM}};
  regs_190 = _RAND_190[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{`RANDOM}};
  regs_191 = _RAND_191[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{`RANDOM}};
  regs_192 = _RAND_192[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{`RANDOM}};
  regs_193 = _RAND_193[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{`RANDOM}};
  regs_194 = _RAND_194[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{`RANDOM}};
  regs_195 = _RAND_195[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{`RANDOM}};
  regs_196 = _RAND_196[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{`RANDOM}};
  regs_197 = _RAND_197[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{`RANDOM}};
  regs_198 = _RAND_198[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{`RANDOM}};
  regs_199 = _RAND_199[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{`RANDOM}};
  regs_200 = _RAND_200[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{`RANDOM}};
  regs_201 = _RAND_201[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{`RANDOM}};
  regs_202 = _RAND_202[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{`RANDOM}};
  regs_203 = _RAND_203[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{`RANDOM}};
  regs_204 = _RAND_204[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{`RANDOM}};
  regs_205 = _RAND_205[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{`RANDOM}};
  regs_206 = _RAND_206[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{`RANDOM}};
  regs_207 = _RAND_207[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{`RANDOM}};
  regs_208 = _RAND_208[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{`RANDOM}};
  regs_209 = _RAND_209[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{`RANDOM}};
  regs_210 = _RAND_210[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{`RANDOM}};
  regs_211 = _RAND_211[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{`RANDOM}};
  regs_212 = _RAND_212[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{`RANDOM}};
  regs_213 = _RAND_213[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{`RANDOM}};
  regs_214 = _RAND_214[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{`RANDOM}};
  regs_215 = _RAND_215[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{`RANDOM}};
  regs_216 = _RAND_216[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{`RANDOM}};
  regs_217 = _RAND_217[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{`RANDOM}};
  regs_218 = _RAND_218[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{`RANDOM}};
  regs_219 = _RAND_219[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{`RANDOM}};
  regs_220 = _RAND_220[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{`RANDOM}};
  regs_221 = _RAND_221[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{`RANDOM}};
  regs_222 = _RAND_222[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{`RANDOM}};
  regs_223 = _RAND_223[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{`RANDOM}};
  regs_224 = _RAND_224[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{`RANDOM}};
  regs_225 = _RAND_225[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{`RANDOM}};
  regs_226 = _RAND_226[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{`RANDOM}};
  regs_227 = _RAND_227[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{`RANDOM}};
  regs_228 = _RAND_228[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{`RANDOM}};
  regs_229 = _RAND_229[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{`RANDOM}};
  regs_230 = _RAND_230[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{`RANDOM}};
  regs_231 = _RAND_231[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{`RANDOM}};
  regs_232 = _RAND_232[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {1{`RANDOM}};
  regs_233 = _RAND_233[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {1{`RANDOM}};
  regs_234 = _RAND_234[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {1{`RANDOM}};
  regs_235 = _RAND_235[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{`RANDOM}};
  regs_236 = _RAND_236[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {1{`RANDOM}};
  regs_237 = _RAND_237[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{`RANDOM}};
  regs_238 = _RAND_238[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {1{`RANDOM}};
  regs_239 = _RAND_239[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{`RANDOM}};
  regs_240 = _RAND_240[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {1{`RANDOM}};
  regs_241 = _RAND_241[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{`RANDOM}};
  regs_242 = _RAND_242[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {1{`RANDOM}};
  regs_243 = _RAND_243[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {1{`RANDOM}};
  regs_244 = _RAND_244[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {1{`RANDOM}};
  regs_245 = _RAND_245[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{`RANDOM}};
  regs_246 = _RAND_246[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {1{`RANDOM}};
  regs_247 = _RAND_247[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {1{`RANDOM}};
  regs_248 = _RAND_248[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {1{`RANDOM}};
  regs_249 = _RAND_249[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {1{`RANDOM}};
  regs_250 = _RAND_250[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_251 = {1{`RANDOM}};
  regs_251 = _RAND_251[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_252 = {1{`RANDOM}};
  regs_252 = _RAND_252[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_253 = {1{`RANDOM}};
  regs_253 = _RAND_253[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_254 = {1{`RANDOM}};
  regs_254 = _RAND_254[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_255 = {1{`RANDOM}};
  regs_255 = _RAND_255[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_256 = {1{`RANDOM}};
  regs_256 = _RAND_256[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_257 = {1{`RANDOM}};
  regs_257 = _RAND_257[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_258 = {1{`RANDOM}};
  regs_258 = _RAND_258[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_259 = {1{`RANDOM}};
  regs_259 = _RAND_259[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_260 = {1{`RANDOM}};
  regs_260 = _RAND_260[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_261 = {1{`RANDOM}};
  regs_261 = _RAND_261[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_262 = {1{`RANDOM}};
  regs_262 = _RAND_262[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_263 = {1{`RANDOM}};
  regs_263 = _RAND_263[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_264 = {1{`RANDOM}};
  regs_264 = _RAND_264[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_265 = {1{`RANDOM}};
  regs_265 = _RAND_265[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_266 = {1{`RANDOM}};
  regs_266 = _RAND_266[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_267 = {1{`RANDOM}};
  regs_267 = _RAND_267[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_268 = {1{`RANDOM}};
  regs_268 = _RAND_268[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_269 = {1{`RANDOM}};
  regs_269 = _RAND_269[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_270 = {1{`RANDOM}};
  regs_270 = _RAND_270[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_271 = {1{`RANDOM}};
  regs_271 = _RAND_271[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_272 = {1{`RANDOM}};
  regs_272 = _RAND_272[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_273 = {1{`RANDOM}};
  regs_273 = _RAND_273[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_274 = {1{`RANDOM}};
  regs_274 = _RAND_274[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_275 = {1{`RANDOM}};
  regs_275 = _RAND_275[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_276 = {1{`RANDOM}};
  regs_276 = _RAND_276[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_277 = {1{`RANDOM}};
  regs_277 = _RAND_277[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_278 = {1{`RANDOM}};
  regs_278 = _RAND_278[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_279 = {1{`RANDOM}};
  regs_279 = _RAND_279[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_280 = {1{`RANDOM}};
  regs_280 = _RAND_280[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_281 = {1{`RANDOM}};
  regs_281 = _RAND_281[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_282 = {1{`RANDOM}};
  regs_282 = _RAND_282[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_283 = {1{`RANDOM}};
  regs_283 = _RAND_283[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_284 = {1{`RANDOM}};
  regs_284 = _RAND_284[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_285 = {1{`RANDOM}};
  regs_285 = _RAND_285[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_286 = {1{`RANDOM}};
  regs_286 = _RAND_286[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_287 = {1{`RANDOM}};
  regs_287 = _RAND_287[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_288 = {1{`RANDOM}};
  regs_288 = _RAND_288[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_289 = {1{`RANDOM}};
  regs_289 = _RAND_289[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_290 = {1{`RANDOM}};
  regs_290 = _RAND_290[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_291 = {1{`RANDOM}};
  regs_291 = _RAND_291[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_292 = {1{`RANDOM}};
  regs_292 = _RAND_292[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_293 = {1{`RANDOM}};
  regs_293 = _RAND_293[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_294 = {1{`RANDOM}};
  regs_294 = _RAND_294[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_295 = {1{`RANDOM}};
  regs_295 = _RAND_295[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_296 = {1{`RANDOM}};
  regs_296 = _RAND_296[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_297 = {1{`RANDOM}};
  regs_297 = _RAND_297[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_298 = {1{`RANDOM}};
  regs_298 = _RAND_298[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_299 = {1{`RANDOM}};
  regs_299 = _RAND_299[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_300 = {1{`RANDOM}};
  regs_300 = _RAND_300[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_301 = {1{`RANDOM}};
  regs_301 = _RAND_301[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_302 = {1{`RANDOM}};
  regs_302 = _RAND_302[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_303 = {1{`RANDOM}};
  regs_303 = _RAND_303[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_304 = {1{`RANDOM}};
  regs_304 = _RAND_304[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_305 = {1{`RANDOM}};
  regs_305 = _RAND_305[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_306 = {1{`RANDOM}};
  regs_306 = _RAND_306[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_307 = {1{`RANDOM}};
  regs_307 = _RAND_307[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_308 = {1{`RANDOM}};
  regs_308 = _RAND_308[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_309 = {1{`RANDOM}};
  regs_309 = _RAND_309[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_310 = {1{`RANDOM}};
  regs_310 = _RAND_310[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_311 = {1{`RANDOM}};
  regs_311 = _RAND_311[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_312 = {1{`RANDOM}};
  regs_312 = _RAND_312[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_313 = {1{`RANDOM}};
  regs_313 = _RAND_313[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_314 = {1{`RANDOM}};
  regs_314 = _RAND_314[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_315 = {1{`RANDOM}};
  regs_315 = _RAND_315[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_316 = {1{`RANDOM}};
  regs_316 = _RAND_316[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_317 = {1{`RANDOM}};
  regs_317 = _RAND_317[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_318 = {1{`RANDOM}};
  regs_318 = _RAND_318[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_319 = {1{`RANDOM}};
  regs_319 = _RAND_319[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_320 = {1{`RANDOM}};
  regs_320 = _RAND_320[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_321 = {1{`RANDOM}};
  regs_321 = _RAND_321[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_322 = {1{`RANDOM}};
  regs_322 = _RAND_322[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_323 = {1{`RANDOM}};
  regs_323 = _RAND_323[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_324 = {1{`RANDOM}};
  regs_324 = _RAND_324[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_325 = {1{`RANDOM}};
  regs_325 = _RAND_325[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_326 = {1{`RANDOM}};
  regs_326 = _RAND_326[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_327 = {1{`RANDOM}};
  regs_327 = _RAND_327[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_328 = {1{`RANDOM}};
  regs_328 = _RAND_328[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_329 = {1{`RANDOM}};
  regs_329 = _RAND_329[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_330 = {1{`RANDOM}};
  regs_330 = _RAND_330[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_331 = {1{`RANDOM}};
  regs_331 = _RAND_331[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_332 = {1{`RANDOM}};
  regs_332 = _RAND_332[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_333 = {1{`RANDOM}};
  regs_333 = _RAND_333[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_334 = {1{`RANDOM}};
  regs_334 = _RAND_334[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_335 = {1{`RANDOM}};
  regs_335 = _RAND_335[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_336 = {1{`RANDOM}};
  regs_336 = _RAND_336[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_337 = {1{`RANDOM}};
  regs_337 = _RAND_337[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_338 = {1{`RANDOM}};
  regs_338 = _RAND_338[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_339 = {1{`RANDOM}};
  regs_339 = _RAND_339[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_340 = {1{`RANDOM}};
  regs_340 = _RAND_340[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_341 = {1{`RANDOM}};
  regs_341 = _RAND_341[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_342 = {1{`RANDOM}};
  regs_342 = _RAND_342[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_343 = {1{`RANDOM}};
  regs_343 = _RAND_343[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_344 = {1{`RANDOM}};
  regs_344 = _RAND_344[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_345 = {1{`RANDOM}};
  regs_345 = _RAND_345[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_346 = {1{`RANDOM}};
  regs_346 = _RAND_346[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_347 = {1{`RANDOM}};
  regs_347 = _RAND_347[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_348 = {1{`RANDOM}};
  regs_348 = _RAND_348[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_349 = {1{`RANDOM}};
  regs_349 = _RAND_349[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_350 = {1{`RANDOM}};
  regs_350 = _RAND_350[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_351 = {1{`RANDOM}};
  regs_351 = _RAND_351[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_352 = {1{`RANDOM}};
  regs_352 = _RAND_352[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_353 = {1{`RANDOM}};
  regs_353 = _RAND_353[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_354 = {1{`RANDOM}};
  regs_354 = _RAND_354[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_355 = {1{`RANDOM}};
  regs_355 = _RAND_355[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_356 = {1{`RANDOM}};
  regs_356 = _RAND_356[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_357 = {1{`RANDOM}};
  regs_357 = _RAND_357[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_358 = {1{`RANDOM}};
  regs_358 = _RAND_358[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_359 = {1{`RANDOM}};
  regs_359 = _RAND_359[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_360 = {1{`RANDOM}};
  regs_360 = _RAND_360[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_361 = {1{`RANDOM}};
  regs_361 = _RAND_361[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_362 = {1{`RANDOM}};
  regs_362 = _RAND_362[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_363 = {1{`RANDOM}};
  regs_363 = _RAND_363[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_364 = {1{`RANDOM}};
  regs_364 = _RAND_364[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_365 = {1{`RANDOM}};
  regs_365 = _RAND_365[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_366 = {1{`RANDOM}};
  regs_366 = _RAND_366[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_367 = {1{`RANDOM}};
  regs_367 = _RAND_367[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_368 = {1{`RANDOM}};
  regs_368 = _RAND_368[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_369 = {1{`RANDOM}};
  regs_369 = _RAND_369[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_370 = {1{`RANDOM}};
  regs_370 = _RAND_370[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_371 = {1{`RANDOM}};
  regs_371 = _RAND_371[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_372 = {1{`RANDOM}};
  regs_372 = _RAND_372[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_373 = {1{`RANDOM}};
  regs_373 = _RAND_373[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_374 = {1{`RANDOM}};
  regs_374 = _RAND_374[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_375 = {1{`RANDOM}};
  regs_375 = _RAND_375[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_376 = {1{`RANDOM}};
  regs_376 = _RAND_376[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_377 = {1{`RANDOM}};
  regs_377 = _RAND_377[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_378 = {1{`RANDOM}};
  regs_378 = _RAND_378[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_379 = {1{`RANDOM}};
  regs_379 = _RAND_379[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_380 = {1{`RANDOM}};
  regs_380 = _RAND_380[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_381 = {1{`RANDOM}};
  regs_381 = _RAND_381[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_382 = {1{`RANDOM}};
  regs_382 = _RAND_382[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_383 = {1{`RANDOM}};
  regs_383 = _RAND_383[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_384 = {1{`RANDOM}};
  regs_384 = _RAND_384[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_385 = {1{`RANDOM}};
  regs_385 = _RAND_385[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_386 = {1{`RANDOM}};
  regs_386 = _RAND_386[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_387 = {1{`RANDOM}};
  regs_387 = _RAND_387[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_388 = {1{`RANDOM}};
  regs_388 = _RAND_388[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_389 = {1{`RANDOM}};
  regs_389 = _RAND_389[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_390 = {1{`RANDOM}};
  regs_390 = _RAND_390[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_391 = {1{`RANDOM}};
  regs_391 = _RAND_391[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_392 = {1{`RANDOM}};
  regs_392 = _RAND_392[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_393 = {1{`RANDOM}};
  regs_393 = _RAND_393[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_394 = {1{`RANDOM}};
  regs_394 = _RAND_394[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_395 = {1{`RANDOM}};
  regs_395 = _RAND_395[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_396 = {1{`RANDOM}};
  regs_396 = _RAND_396[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_397 = {1{`RANDOM}};
  regs_397 = _RAND_397[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_398 = {1{`RANDOM}};
  regs_398 = _RAND_398[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_399 = {1{`RANDOM}};
  regs_399 = _RAND_399[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      regs_0 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_0 <= io_in_bits;
      end
    end
    if (reset) begin
      regs_1 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_1 <= regs_0;
      end
    end
    if (reset) begin
      regs_2 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_2 <= regs_1;
      end
    end
    if (reset) begin
      regs_3 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_3 <= regs_2;
      end
    end
    if (reset) begin
      regs_4 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_4 <= regs_3;
      end
    end
    if (reset) begin
      regs_5 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_5 <= regs_4;
      end
    end
    if (reset) begin
      regs_6 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_6 <= regs_5;
      end
    end
    if (reset) begin
      regs_7 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_7 <= regs_6;
      end
    end
    if (reset) begin
      regs_8 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_8 <= regs_7;
      end
    end
    if (reset) begin
      regs_9 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_9 <= regs_8;
      end
    end
    if (reset) begin
      regs_10 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_10 <= regs_9;
      end
    end
    if (reset) begin
      regs_11 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_11 <= regs_10;
      end
    end
    if (reset) begin
      regs_12 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_12 <= regs_11;
      end
    end
    if (reset) begin
      regs_13 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_13 <= regs_12;
      end
    end
    if (reset) begin
      regs_14 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_14 <= regs_13;
      end
    end
    if (reset) begin
      regs_15 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_15 <= regs_14;
      end
    end
    if (reset) begin
      regs_16 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_16 <= regs_15;
      end
    end
    if (reset) begin
      regs_17 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_17 <= regs_16;
      end
    end
    if (reset) begin
      regs_18 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_18 <= regs_17;
      end
    end
    if (reset) begin
      regs_19 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_19 <= regs_18;
      end
    end
    if (reset) begin
      regs_20 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_20 <= regs_19;
      end
    end
    if (reset) begin
      regs_21 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_21 <= regs_20;
      end
    end
    if (reset) begin
      regs_22 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_22 <= regs_21;
      end
    end
    if (reset) begin
      regs_23 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_23 <= regs_22;
      end
    end
    if (reset) begin
      regs_24 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_24 <= regs_23;
      end
    end
    if (reset) begin
      regs_25 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_25 <= regs_24;
      end
    end
    if (reset) begin
      regs_26 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_26 <= regs_25;
      end
    end
    if (reset) begin
      regs_27 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_27 <= regs_26;
      end
    end
    if (reset) begin
      regs_28 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_28 <= regs_27;
      end
    end
    if (reset) begin
      regs_29 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_29 <= regs_28;
      end
    end
    if (reset) begin
      regs_30 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_30 <= regs_29;
      end
    end
    if (reset) begin
      regs_31 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_31 <= regs_30;
      end
    end
    if (reset) begin
      regs_32 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_32 <= regs_31;
      end
    end
    if (reset) begin
      regs_33 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_33 <= regs_32;
      end
    end
    if (reset) begin
      regs_34 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_34 <= regs_33;
      end
    end
    if (reset) begin
      regs_35 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_35 <= regs_34;
      end
    end
    if (reset) begin
      regs_36 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_36 <= regs_35;
      end
    end
    if (reset) begin
      regs_37 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_37 <= regs_36;
      end
    end
    if (reset) begin
      regs_38 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_38 <= regs_37;
      end
    end
    if (reset) begin
      regs_39 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_39 <= regs_38;
      end
    end
    if (reset) begin
      regs_40 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_40 <= regs_39;
      end
    end
    if (reset) begin
      regs_41 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_41 <= regs_40;
      end
    end
    if (reset) begin
      regs_42 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_42 <= regs_41;
      end
    end
    if (reset) begin
      regs_43 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_43 <= regs_42;
      end
    end
    if (reset) begin
      regs_44 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_44 <= regs_43;
      end
    end
    if (reset) begin
      regs_45 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_45 <= regs_44;
      end
    end
    if (reset) begin
      regs_46 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_46 <= regs_45;
      end
    end
    if (reset) begin
      regs_47 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_47 <= regs_46;
      end
    end
    if (reset) begin
      regs_48 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_48 <= regs_47;
      end
    end
    if (reset) begin
      regs_49 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_49 <= regs_48;
      end
    end
    if (reset) begin
      regs_50 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_50 <= regs_49;
      end
    end
    if (reset) begin
      regs_51 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_51 <= regs_50;
      end
    end
    if (reset) begin
      regs_52 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_52 <= regs_51;
      end
    end
    if (reset) begin
      regs_53 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_53 <= regs_52;
      end
    end
    if (reset) begin
      regs_54 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_54 <= regs_53;
      end
    end
    if (reset) begin
      regs_55 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_55 <= regs_54;
      end
    end
    if (reset) begin
      regs_56 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_56 <= regs_55;
      end
    end
    if (reset) begin
      regs_57 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_57 <= regs_56;
      end
    end
    if (reset) begin
      regs_58 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_58 <= regs_57;
      end
    end
    if (reset) begin
      regs_59 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_59 <= regs_58;
      end
    end
    if (reset) begin
      regs_60 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_60 <= regs_59;
      end
    end
    if (reset) begin
      regs_61 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_61 <= regs_60;
      end
    end
    if (reset) begin
      regs_62 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_62 <= regs_61;
      end
    end
    if (reset) begin
      regs_63 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_63 <= regs_62;
      end
    end
    if (reset) begin
      regs_64 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_64 <= regs_63;
      end
    end
    if (reset) begin
      regs_65 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_65 <= regs_64;
      end
    end
    if (reset) begin
      regs_66 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_66 <= regs_65;
      end
    end
    if (reset) begin
      regs_67 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_67 <= regs_66;
      end
    end
    if (reset) begin
      regs_68 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_68 <= regs_67;
      end
    end
    if (reset) begin
      regs_69 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_69 <= regs_68;
      end
    end
    if (reset) begin
      regs_70 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_70 <= regs_69;
      end
    end
    if (reset) begin
      regs_71 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_71 <= regs_70;
      end
    end
    if (reset) begin
      regs_72 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_72 <= regs_71;
      end
    end
    if (reset) begin
      regs_73 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_73 <= regs_72;
      end
    end
    if (reset) begin
      regs_74 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_74 <= regs_73;
      end
    end
    if (reset) begin
      regs_75 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_75 <= regs_74;
      end
    end
    if (reset) begin
      regs_76 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_76 <= regs_75;
      end
    end
    if (reset) begin
      regs_77 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_77 <= regs_76;
      end
    end
    if (reset) begin
      regs_78 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_78 <= regs_77;
      end
    end
    if (reset) begin
      regs_79 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_79 <= regs_78;
      end
    end
    if (reset) begin
      regs_80 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_80 <= regs_79;
      end
    end
    if (reset) begin
      regs_81 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_81 <= regs_80;
      end
    end
    if (reset) begin
      regs_82 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_82 <= regs_81;
      end
    end
    if (reset) begin
      regs_83 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_83 <= regs_82;
      end
    end
    if (reset) begin
      regs_84 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_84 <= regs_83;
      end
    end
    if (reset) begin
      regs_85 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_85 <= regs_84;
      end
    end
    if (reset) begin
      regs_86 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_86 <= regs_85;
      end
    end
    if (reset) begin
      regs_87 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_87 <= regs_86;
      end
    end
    if (reset) begin
      regs_88 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_88 <= regs_87;
      end
    end
    if (reset) begin
      regs_89 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_89 <= regs_88;
      end
    end
    if (reset) begin
      regs_90 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_90 <= regs_89;
      end
    end
    if (reset) begin
      regs_91 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_91 <= regs_90;
      end
    end
    if (reset) begin
      regs_92 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_92 <= regs_91;
      end
    end
    if (reset) begin
      regs_93 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_93 <= regs_92;
      end
    end
    if (reset) begin
      regs_94 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_94 <= regs_93;
      end
    end
    if (reset) begin
      regs_95 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_95 <= regs_94;
      end
    end
    if (reset) begin
      regs_96 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_96 <= regs_95;
      end
    end
    if (reset) begin
      regs_97 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_97 <= regs_96;
      end
    end
    if (reset) begin
      regs_98 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_98 <= regs_97;
      end
    end
    if (reset) begin
      regs_99 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_99 <= regs_98;
      end
    end
    if (reset) begin
      regs_100 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_100 <= regs_99;
      end
    end
    if (reset) begin
      regs_101 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_101 <= regs_100;
      end
    end
    if (reset) begin
      regs_102 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_102 <= regs_101;
      end
    end
    if (reset) begin
      regs_103 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_103 <= regs_102;
      end
    end
    if (reset) begin
      regs_104 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_104 <= regs_103;
      end
    end
    if (reset) begin
      regs_105 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_105 <= regs_104;
      end
    end
    if (reset) begin
      regs_106 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_106 <= regs_105;
      end
    end
    if (reset) begin
      regs_107 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_107 <= regs_106;
      end
    end
    if (reset) begin
      regs_108 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_108 <= regs_107;
      end
    end
    if (reset) begin
      regs_109 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_109 <= regs_108;
      end
    end
    if (reset) begin
      regs_110 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_110 <= regs_109;
      end
    end
    if (reset) begin
      regs_111 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_111 <= regs_110;
      end
    end
    if (reset) begin
      regs_112 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_112 <= regs_111;
      end
    end
    if (reset) begin
      regs_113 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_113 <= regs_112;
      end
    end
    if (reset) begin
      regs_114 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_114 <= regs_113;
      end
    end
    if (reset) begin
      regs_115 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_115 <= regs_114;
      end
    end
    if (reset) begin
      regs_116 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_116 <= regs_115;
      end
    end
    if (reset) begin
      regs_117 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_117 <= regs_116;
      end
    end
    if (reset) begin
      regs_118 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_118 <= regs_117;
      end
    end
    if (reset) begin
      regs_119 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_119 <= regs_118;
      end
    end
    if (reset) begin
      regs_120 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_120 <= regs_119;
      end
    end
    if (reset) begin
      regs_121 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_121 <= regs_120;
      end
    end
    if (reset) begin
      regs_122 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_122 <= regs_121;
      end
    end
    if (reset) begin
      regs_123 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_123 <= regs_122;
      end
    end
    if (reset) begin
      regs_124 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_124 <= regs_123;
      end
    end
    if (reset) begin
      regs_125 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_125 <= regs_124;
      end
    end
    if (reset) begin
      regs_126 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_126 <= regs_125;
      end
    end
    if (reset) begin
      regs_127 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_127 <= regs_126;
      end
    end
    if (reset) begin
      regs_128 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_128 <= regs_127;
      end
    end
    if (reset) begin
      regs_129 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_129 <= regs_128;
      end
    end
    if (reset) begin
      regs_130 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_130 <= regs_129;
      end
    end
    if (reset) begin
      regs_131 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_131 <= regs_130;
      end
    end
    if (reset) begin
      regs_132 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_132 <= regs_131;
      end
    end
    if (reset) begin
      regs_133 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_133 <= regs_132;
      end
    end
    if (reset) begin
      regs_134 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_134 <= regs_133;
      end
    end
    if (reset) begin
      regs_135 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_135 <= regs_134;
      end
    end
    if (reset) begin
      regs_136 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_136 <= regs_135;
      end
    end
    if (reset) begin
      regs_137 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_137 <= regs_136;
      end
    end
    if (reset) begin
      regs_138 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_138 <= regs_137;
      end
    end
    if (reset) begin
      regs_139 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_139 <= regs_138;
      end
    end
    if (reset) begin
      regs_140 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_140 <= regs_139;
      end
    end
    if (reset) begin
      regs_141 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_141 <= regs_140;
      end
    end
    if (reset) begin
      regs_142 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_142 <= regs_141;
      end
    end
    if (reset) begin
      regs_143 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_143 <= regs_142;
      end
    end
    if (reset) begin
      regs_144 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_144 <= regs_143;
      end
    end
    if (reset) begin
      regs_145 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_145 <= regs_144;
      end
    end
    if (reset) begin
      regs_146 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_146 <= regs_145;
      end
    end
    if (reset) begin
      regs_147 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_147 <= regs_146;
      end
    end
    if (reset) begin
      regs_148 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_148 <= regs_147;
      end
    end
    if (reset) begin
      regs_149 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_149 <= regs_148;
      end
    end
    if (reset) begin
      regs_150 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_150 <= regs_149;
      end
    end
    if (reset) begin
      regs_151 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_151 <= regs_150;
      end
    end
    if (reset) begin
      regs_152 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_152 <= regs_151;
      end
    end
    if (reset) begin
      regs_153 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_153 <= regs_152;
      end
    end
    if (reset) begin
      regs_154 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_154 <= regs_153;
      end
    end
    if (reset) begin
      regs_155 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_155 <= regs_154;
      end
    end
    if (reset) begin
      regs_156 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_156 <= regs_155;
      end
    end
    if (reset) begin
      regs_157 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_157 <= regs_156;
      end
    end
    if (reset) begin
      regs_158 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_158 <= regs_157;
      end
    end
    if (reset) begin
      regs_159 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_159 <= regs_158;
      end
    end
    if (reset) begin
      regs_160 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_160 <= regs_159;
      end
    end
    if (reset) begin
      regs_161 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_161 <= regs_160;
      end
    end
    if (reset) begin
      regs_162 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_162 <= regs_161;
      end
    end
    if (reset) begin
      regs_163 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_163 <= regs_162;
      end
    end
    if (reset) begin
      regs_164 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_164 <= regs_163;
      end
    end
    if (reset) begin
      regs_165 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_165 <= regs_164;
      end
    end
    if (reset) begin
      regs_166 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_166 <= regs_165;
      end
    end
    if (reset) begin
      regs_167 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_167 <= regs_166;
      end
    end
    if (reset) begin
      regs_168 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_168 <= regs_167;
      end
    end
    if (reset) begin
      regs_169 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_169 <= regs_168;
      end
    end
    if (reset) begin
      regs_170 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_170 <= regs_169;
      end
    end
    if (reset) begin
      regs_171 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_171 <= regs_170;
      end
    end
    if (reset) begin
      regs_172 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_172 <= regs_171;
      end
    end
    if (reset) begin
      regs_173 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_173 <= regs_172;
      end
    end
    if (reset) begin
      regs_174 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_174 <= regs_173;
      end
    end
    if (reset) begin
      regs_175 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_175 <= regs_174;
      end
    end
    if (reset) begin
      regs_176 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_176 <= regs_175;
      end
    end
    if (reset) begin
      regs_177 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_177 <= regs_176;
      end
    end
    if (reset) begin
      regs_178 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_178 <= regs_177;
      end
    end
    if (reset) begin
      regs_179 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_179 <= regs_178;
      end
    end
    if (reset) begin
      regs_180 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_180 <= regs_179;
      end
    end
    if (reset) begin
      regs_181 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_181 <= regs_180;
      end
    end
    if (reset) begin
      regs_182 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_182 <= regs_181;
      end
    end
    if (reset) begin
      regs_183 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_183 <= regs_182;
      end
    end
    if (reset) begin
      regs_184 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_184 <= regs_183;
      end
    end
    if (reset) begin
      regs_185 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_185 <= regs_184;
      end
    end
    if (reset) begin
      regs_186 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_186 <= regs_185;
      end
    end
    if (reset) begin
      regs_187 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_187 <= regs_186;
      end
    end
    if (reset) begin
      regs_188 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_188 <= regs_187;
      end
    end
    if (reset) begin
      regs_189 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_189 <= regs_188;
      end
    end
    if (reset) begin
      regs_190 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_190 <= regs_189;
      end
    end
    if (reset) begin
      regs_191 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_191 <= regs_190;
      end
    end
    if (reset) begin
      regs_192 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_192 <= regs_191;
      end
    end
    if (reset) begin
      regs_193 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_193 <= regs_192;
      end
    end
    if (reset) begin
      regs_194 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_194 <= regs_193;
      end
    end
    if (reset) begin
      regs_195 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_195 <= regs_194;
      end
    end
    if (reset) begin
      regs_196 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_196 <= regs_195;
      end
    end
    if (reset) begin
      regs_197 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_197 <= regs_196;
      end
    end
    if (reset) begin
      regs_198 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_198 <= regs_197;
      end
    end
    if (reset) begin
      regs_199 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_199 <= regs_198;
      end
    end
    if (reset) begin
      regs_200 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_200 <= regs_199;
      end
    end
    if (reset) begin
      regs_201 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_201 <= regs_200;
      end
    end
    if (reset) begin
      regs_202 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_202 <= regs_201;
      end
    end
    if (reset) begin
      regs_203 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_203 <= regs_202;
      end
    end
    if (reset) begin
      regs_204 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_204 <= regs_203;
      end
    end
    if (reset) begin
      regs_205 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_205 <= regs_204;
      end
    end
    if (reset) begin
      regs_206 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_206 <= regs_205;
      end
    end
    if (reset) begin
      regs_207 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_207 <= regs_206;
      end
    end
    if (reset) begin
      regs_208 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_208 <= regs_207;
      end
    end
    if (reset) begin
      regs_209 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_209 <= regs_208;
      end
    end
    if (reset) begin
      regs_210 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_210 <= regs_209;
      end
    end
    if (reset) begin
      regs_211 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_211 <= regs_210;
      end
    end
    if (reset) begin
      regs_212 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_212 <= regs_211;
      end
    end
    if (reset) begin
      regs_213 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_213 <= regs_212;
      end
    end
    if (reset) begin
      regs_214 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_214 <= regs_213;
      end
    end
    if (reset) begin
      regs_215 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_215 <= regs_214;
      end
    end
    if (reset) begin
      regs_216 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_216 <= regs_215;
      end
    end
    if (reset) begin
      regs_217 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_217 <= regs_216;
      end
    end
    if (reset) begin
      regs_218 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_218 <= regs_217;
      end
    end
    if (reset) begin
      regs_219 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_219 <= regs_218;
      end
    end
    if (reset) begin
      regs_220 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_220 <= regs_219;
      end
    end
    if (reset) begin
      regs_221 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_221 <= regs_220;
      end
    end
    if (reset) begin
      regs_222 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_222 <= regs_221;
      end
    end
    if (reset) begin
      regs_223 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_223 <= regs_222;
      end
    end
    if (reset) begin
      regs_224 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_224 <= regs_223;
      end
    end
    if (reset) begin
      regs_225 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_225 <= regs_224;
      end
    end
    if (reset) begin
      regs_226 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_226 <= regs_225;
      end
    end
    if (reset) begin
      regs_227 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_227 <= regs_226;
      end
    end
    if (reset) begin
      regs_228 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_228 <= regs_227;
      end
    end
    if (reset) begin
      regs_229 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_229 <= regs_228;
      end
    end
    if (reset) begin
      regs_230 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_230 <= regs_229;
      end
    end
    if (reset) begin
      regs_231 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_231 <= regs_230;
      end
    end
    if (reset) begin
      regs_232 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_232 <= regs_231;
      end
    end
    if (reset) begin
      regs_233 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_233 <= regs_232;
      end
    end
    if (reset) begin
      regs_234 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_234 <= regs_233;
      end
    end
    if (reset) begin
      regs_235 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_235 <= regs_234;
      end
    end
    if (reset) begin
      regs_236 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_236 <= regs_235;
      end
    end
    if (reset) begin
      regs_237 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_237 <= regs_236;
      end
    end
    if (reset) begin
      regs_238 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_238 <= regs_237;
      end
    end
    if (reset) begin
      regs_239 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_239 <= regs_238;
      end
    end
    if (reset) begin
      regs_240 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_240 <= regs_239;
      end
    end
    if (reset) begin
      regs_241 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_241 <= regs_240;
      end
    end
    if (reset) begin
      regs_242 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_242 <= regs_241;
      end
    end
    if (reset) begin
      regs_243 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_243 <= regs_242;
      end
    end
    if (reset) begin
      regs_244 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_244 <= regs_243;
      end
    end
    if (reset) begin
      regs_245 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_245 <= regs_244;
      end
    end
    if (reset) begin
      regs_246 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_246 <= regs_245;
      end
    end
    if (reset) begin
      regs_247 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_247 <= regs_246;
      end
    end
    if (reset) begin
      regs_248 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_248 <= regs_247;
      end
    end
    if (reset) begin
      regs_249 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_249 <= regs_248;
      end
    end
    if (reset) begin
      regs_250 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_250 <= regs_249;
      end
    end
    if (reset) begin
      regs_251 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_251 <= regs_250;
      end
    end
    if (reset) begin
      regs_252 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_252 <= regs_251;
      end
    end
    if (reset) begin
      regs_253 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_253 <= regs_252;
      end
    end
    if (reset) begin
      regs_254 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_254 <= regs_253;
      end
    end
    if (reset) begin
      regs_255 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_255 <= regs_254;
      end
    end
    if (reset) begin
      regs_256 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_256 <= regs_255;
      end
    end
    if (reset) begin
      regs_257 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_257 <= regs_256;
      end
    end
    if (reset) begin
      regs_258 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_258 <= regs_257;
      end
    end
    if (reset) begin
      regs_259 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_259 <= regs_258;
      end
    end
    if (reset) begin
      regs_260 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_260 <= regs_259;
      end
    end
    if (reset) begin
      regs_261 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_261 <= regs_260;
      end
    end
    if (reset) begin
      regs_262 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_262 <= regs_261;
      end
    end
    if (reset) begin
      regs_263 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_263 <= regs_262;
      end
    end
    if (reset) begin
      regs_264 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_264 <= regs_263;
      end
    end
    if (reset) begin
      regs_265 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_265 <= regs_264;
      end
    end
    if (reset) begin
      regs_266 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_266 <= regs_265;
      end
    end
    if (reset) begin
      regs_267 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_267 <= regs_266;
      end
    end
    if (reset) begin
      regs_268 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_268 <= regs_267;
      end
    end
    if (reset) begin
      regs_269 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_269 <= regs_268;
      end
    end
    if (reset) begin
      regs_270 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_270 <= regs_269;
      end
    end
    if (reset) begin
      regs_271 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_271 <= regs_270;
      end
    end
    if (reset) begin
      regs_272 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_272 <= regs_271;
      end
    end
    if (reset) begin
      regs_273 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_273 <= regs_272;
      end
    end
    if (reset) begin
      regs_274 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_274 <= regs_273;
      end
    end
    if (reset) begin
      regs_275 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_275 <= regs_274;
      end
    end
    if (reset) begin
      regs_276 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_276 <= regs_275;
      end
    end
    if (reset) begin
      regs_277 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_277 <= regs_276;
      end
    end
    if (reset) begin
      regs_278 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_278 <= regs_277;
      end
    end
    if (reset) begin
      regs_279 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_279 <= regs_278;
      end
    end
    if (reset) begin
      regs_280 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_280 <= regs_279;
      end
    end
    if (reset) begin
      regs_281 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_281 <= regs_280;
      end
    end
    if (reset) begin
      regs_282 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_282 <= regs_281;
      end
    end
    if (reset) begin
      regs_283 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_283 <= regs_282;
      end
    end
    if (reset) begin
      regs_284 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_284 <= regs_283;
      end
    end
    if (reset) begin
      regs_285 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_285 <= regs_284;
      end
    end
    if (reset) begin
      regs_286 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_286 <= regs_285;
      end
    end
    if (reset) begin
      regs_287 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_287 <= regs_286;
      end
    end
    if (reset) begin
      regs_288 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_288 <= regs_287;
      end
    end
    if (reset) begin
      regs_289 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_289 <= regs_288;
      end
    end
    if (reset) begin
      regs_290 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_290 <= regs_289;
      end
    end
    if (reset) begin
      regs_291 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_291 <= regs_290;
      end
    end
    if (reset) begin
      regs_292 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_292 <= regs_291;
      end
    end
    if (reset) begin
      regs_293 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_293 <= regs_292;
      end
    end
    if (reset) begin
      regs_294 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_294 <= regs_293;
      end
    end
    if (reset) begin
      regs_295 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_295 <= regs_294;
      end
    end
    if (reset) begin
      regs_296 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_296 <= regs_295;
      end
    end
    if (reset) begin
      regs_297 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_297 <= regs_296;
      end
    end
    if (reset) begin
      regs_298 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_298 <= regs_297;
      end
    end
    if (reset) begin
      regs_299 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_299 <= regs_298;
      end
    end
    if (reset) begin
      regs_300 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_300 <= regs_299;
      end
    end
    if (reset) begin
      regs_301 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_301 <= regs_300;
      end
    end
    if (reset) begin
      regs_302 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_302 <= regs_301;
      end
    end
    if (reset) begin
      regs_303 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_303 <= regs_302;
      end
    end
    if (reset) begin
      regs_304 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_304 <= regs_303;
      end
    end
    if (reset) begin
      regs_305 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_305 <= regs_304;
      end
    end
    if (reset) begin
      regs_306 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_306 <= regs_305;
      end
    end
    if (reset) begin
      regs_307 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_307 <= regs_306;
      end
    end
    if (reset) begin
      regs_308 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_308 <= regs_307;
      end
    end
    if (reset) begin
      regs_309 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_309 <= regs_308;
      end
    end
    if (reset) begin
      regs_310 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_310 <= regs_309;
      end
    end
    if (reset) begin
      regs_311 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_311 <= regs_310;
      end
    end
    if (reset) begin
      regs_312 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_312 <= regs_311;
      end
    end
    if (reset) begin
      regs_313 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_313 <= regs_312;
      end
    end
    if (reset) begin
      regs_314 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_314 <= regs_313;
      end
    end
    if (reset) begin
      regs_315 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_315 <= regs_314;
      end
    end
    if (reset) begin
      regs_316 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_316 <= regs_315;
      end
    end
    if (reset) begin
      regs_317 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_317 <= regs_316;
      end
    end
    if (reset) begin
      regs_318 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_318 <= regs_317;
      end
    end
    if (reset) begin
      regs_319 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_319 <= regs_318;
      end
    end
    if (reset) begin
      regs_320 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_320 <= regs_319;
      end
    end
    if (reset) begin
      regs_321 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_321 <= regs_320;
      end
    end
    if (reset) begin
      regs_322 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_322 <= regs_321;
      end
    end
    if (reset) begin
      regs_323 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_323 <= regs_322;
      end
    end
    if (reset) begin
      regs_324 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_324 <= regs_323;
      end
    end
    if (reset) begin
      regs_325 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_325 <= regs_324;
      end
    end
    if (reset) begin
      regs_326 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_326 <= regs_325;
      end
    end
    if (reset) begin
      regs_327 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_327 <= regs_326;
      end
    end
    if (reset) begin
      regs_328 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_328 <= regs_327;
      end
    end
    if (reset) begin
      regs_329 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_329 <= regs_328;
      end
    end
    if (reset) begin
      regs_330 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_330 <= regs_329;
      end
    end
    if (reset) begin
      regs_331 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_331 <= regs_330;
      end
    end
    if (reset) begin
      regs_332 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_332 <= regs_331;
      end
    end
    if (reset) begin
      regs_333 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_333 <= regs_332;
      end
    end
    if (reset) begin
      regs_334 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_334 <= regs_333;
      end
    end
    if (reset) begin
      regs_335 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_335 <= regs_334;
      end
    end
    if (reset) begin
      regs_336 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_336 <= regs_335;
      end
    end
    if (reset) begin
      regs_337 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_337 <= regs_336;
      end
    end
    if (reset) begin
      regs_338 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_338 <= regs_337;
      end
    end
    if (reset) begin
      regs_339 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_339 <= regs_338;
      end
    end
    if (reset) begin
      regs_340 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_340 <= regs_339;
      end
    end
    if (reset) begin
      regs_341 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_341 <= regs_340;
      end
    end
    if (reset) begin
      regs_342 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_342 <= regs_341;
      end
    end
    if (reset) begin
      regs_343 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_343 <= regs_342;
      end
    end
    if (reset) begin
      regs_344 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_344 <= regs_343;
      end
    end
    if (reset) begin
      regs_345 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_345 <= regs_344;
      end
    end
    if (reset) begin
      regs_346 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_346 <= regs_345;
      end
    end
    if (reset) begin
      regs_347 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_347 <= regs_346;
      end
    end
    if (reset) begin
      regs_348 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_348 <= regs_347;
      end
    end
    if (reset) begin
      regs_349 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_349 <= regs_348;
      end
    end
    if (reset) begin
      regs_350 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_350 <= regs_349;
      end
    end
    if (reset) begin
      regs_351 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_351 <= regs_350;
      end
    end
    if (reset) begin
      regs_352 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_352 <= regs_351;
      end
    end
    if (reset) begin
      regs_353 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_353 <= regs_352;
      end
    end
    if (reset) begin
      regs_354 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_354 <= regs_353;
      end
    end
    if (reset) begin
      regs_355 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_355 <= regs_354;
      end
    end
    if (reset) begin
      regs_356 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_356 <= regs_355;
      end
    end
    if (reset) begin
      regs_357 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_357 <= regs_356;
      end
    end
    if (reset) begin
      regs_358 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_358 <= regs_357;
      end
    end
    if (reset) begin
      regs_359 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_359 <= regs_358;
      end
    end
    if (reset) begin
      regs_360 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_360 <= regs_359;
      end
    end
    if (reset) begin
      regs_361 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_361 <= regs_360;
      end
    end
    if (reset) begin
      regs_362 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_362 <= regs_361;
      end
    end
    if (reset) begin
      regs_363 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_363 <= regs_362;
      end
    end
    if (reset) begin
      regs_364 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_364 <= regs_363;
      end
    end
    if (reset) begin
      regs_365 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_365 <= regs_364;
      end
    end
    if (reset) begin
      regs_366 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_366 <= regs_365;
      end
    end
    if (reset) begin
      regs_367 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_367 <= regs_366;
      end
    end
    if (reset) begin
      regs_368 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_368 <= regs_367;
      end
    end
    if (reset) begin
      regs_369 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_369 <= regs_368;
      end
    end
    if (reset) begin
      regs_370 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_370 <= regs_369;
      end
    end
    if (reset) begin
      regs_371 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_371 <= regs_370;
      end
    end
    if (reset) begin
      regs_372 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_372 <= regs_371;
      end
    end
    if (reset) begin
      regs_373 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_373 <= regs_372;
      end
    end
    if (reset) begin
      regs_374 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_374 <= regs_373;
      end
    end
    if (reset) begin
      regs_375 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_375 <= regs_374;
      end
    end
    if (reset) begin
      regs_376 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_376 <= regs_375;
      end
    end
    if (reset) begin
      regs_377 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_377 <= regs_376;
      end
    end
    if (reset) begin
      regs_378 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_378 <= regs_377;
      end
    end
    if (reset) begin
      regs_379 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_379 <= regs_378;
      end
    end
    if (reset) begin
      regs_380 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_380 <= regs_379;
      end
    end
    if (reset) begin
      regs_381 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_381 <= regs_380;
      end
    end
    if (reset) begin
      regs_382 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_382 <= regs_381;
      end
    end
    if (reset) begin
      regs_383 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_383 <= regs_382;
      end
    end
    if (reset) begin
      regs_384 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_384 <= regs_383;
      end
    end
    if (reset) begin
      regs_385 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_385 <= regs_384;
      end
    end
    if (reset) begin
      regs_386 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_386 <= regs_385;
      end
    end
    if (reset) begin
      regs_387 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_387 <= regs_386;
      end
    end
    if (reset) begin
      regs_388 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_388 <= regs_387;
      end
    end
    if (reset) begin
      regs_389 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_389 <= regs_388;
      end
    end
    if (reset) begin
      regs_390 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_390 <= regs_389;
      end
    end
    if (reset) begin
      regs_391 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_391 <= regs_390;
      end
    end
    if (reset) begin
      regs_392 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_392 <= regs_391;
      end
    end
    if (reset) begin
      regs_393 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_393 <= regs_392;
      end
    end
    if (reset) begin
      regs_394 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_394 <= regs_393;
      end
    end
    if (reset) begin
      regs_395 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_395 <= regs_394;
      end
    end
    if (reset) begin
      regs_396 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_396 <= regs_395;
      end
    end
    if (reset) begin
      regs_397 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_397 <= regs_396;
      end
    end
    if (reset) begin
      regs_398 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_398 <= regs_397;
      end
    end
    if (reset) begin
      regs_399 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_399 <= regs_398;
      end
    end
  end
endmodule
module MemoryBuffer_1(
  input         clock,
  input         reset,
  input         io_in_valid,
  input  [31:0] io_in_bits,
  output [31:0] io_out_bits_0_0,
  output [31:0] io_out_bits_0_1,
  output [31:0] io_out_bits_0_2,
  output [31:0] io_out_bits_0_3,
  output [31:0] io_out_bits_0_4,
  output [31:0] io_out_bits_0_5,
  output [31:0] io_out_bits_0_6,
  output [31:0] io_out_bits_0_7,
  output [31:0] io_out_bits_0_8,
  output [31:0] io_out_bits_0_9,
  output [31:0] io_out_bits_0_10,
  output [31:0] io_out_bits_0_11,
  output [31:0] io_out_bits_0_12,
  output [31:0] io_out_bits_0_13,
  output [31:0] io_out_bits_0_14,
  output [31:0] io_out_bits_0_15,
  output [31:0] io_out_bits_0_16,
  output [31:0] io_out_bits_0_17,
  output [31:0] io_out_bits_0_18,
  output [31:0] io_out_bits_0_19,
  output [31:0] io_out_bits_0_20,
  output [31:0] io_out_bits_0_21,
  output [31:0] io_out_bits_0_22,
  output [31:0] io_out_bits_0_23,
  output [31:0] io_out_bits_0_24,
  output [31:0] io_out_bits_0_25,
  output [31:0] io_out_bits_0_26,
  output [31:0] io_out_bits_0_27,
  output [31:0] io_out_bits_0_28,
  output [31:0] io_out_bits_0_29,
  output [31:0] io_out_bits_0_30,
  output [31:0] io_out_bits_0_31,
  output [31:0] io_out_bits_0_32,
  output [31:0] io_out_bits_0_33,
  output [31:0] io_out_bits_0_34,
  output [31:0] io_out_bits_0_35,
  output [31:0] io_out_bits_0_36,
  output [31:0] io_out_bits_0_37,
  output [31:0] io_out_bits_0_38,
  output [31:0] io_out_bits_0_39,
  output [31:0] io_out_bits_0_40,
  output [31:0] io_out_bits_0_41,
  output [31:0] io_out_bits_0_42,
  output [31:0] io_out_bits_0_43,
  output [31:0] io_out_bits_0_44,
  output [31:0] io_out_bits_0_45,
  output [31:0] io_out_bits_0_46,
  output [31:0] io_out_bits_0_47,
  output [31:0] io_out_bits_0_48,
  output [31:0] io_out_bits_0_49,
  output [31:0] io_out_bits_0_50,
  output [31:0] io_out_bits_0_51,
  output [31:0] io_out_bits_0_52,
  output [31:0] io_out_bits_0_53,
  output [31:0] io_out_bits_0_54,
  output [31:0] io_out_bits_0_55,
  output [31:0] io_out_bits_0_56,
  output [31:0] io_out_bits_0_57,
  output [31:0] io_out_bits_0_58,
  output [31:0] io_out_bits_0_59,
  output [31:0] io_out_bits_0_60,
  output [31:0] io_out_bits_0_61,
  output [31:0] io_out_bits_0_62,
  output [31:0] io_out_bits_0_63,
  output [31:0] io_out_bits_0_64,
  output [31:0] io_out_bits_0_65,
  output [31:0] io_out_bits_0_66,
  output [31:0] io_out_bits_0_67,
  output [31:0] io_out_bits_0_68,
  output [31:0] io_out_bits_0_69,
  output [31:0] io_out_bits_0_70,
  output [31:0] io_out_bits_0_71,
  output [31:0] io_out_bits_0_72,
  output [31:0] io_out_bits_0_73,
  output [31:0] io_out_bits_0_74,
  output [31:0] io_out_bits_0_75,
  output [31:0] io_out_bits_0_76,
  output [31:0] io_out_bits_0_77,
  output [31:0] io_out_bits_0_78,
  output [31:0] io_out_bits_0_79,
  output [31:0] io_out_bits_0_80,
  output [31:0] io_out_bits_0_81,
  output [31:0] io_out_bits_0_82,
  output [31:0] io_out_bits_0_83,
  output [31:0] io_out_bits_0_84,
  output [31:0] io_out_bits_0_85,
  output [31:0] io_out_bits_0_86,
  output [31:0] io_out_bits_0_87,
  output [31:0] io_out_bits_0_88,
  output [31:0] io_out_bits_0_89,
  output [31:0] io_out_bits_0_90,
  output [31:0] io_out_bits_0_91,
  output [31:0] io_out_bits_0_92,
  output [31:0] io_out_bits_0_93,
  output [31:0] io_out_bits_0_94,
  output [31:0] io_out_bits_0_95,
  output [31:0] io_out_bits_0_96,
  output [31:0] io_out_bits_0_97,
  output [31:0] io_out_bits_0_98,
  output [31:0] io_out_bits_0_99
);
  reg [31:0] regs_0; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_0;
  reg [31:0] regs_1; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_1;
  reg [31:0] regs_2; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_2;
  reg [31:0] regs_3; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_3;
  reg [31:0] regs_4; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_4;
  reg [31:0] regs_5; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_5;
  reg [31:0] regs_6; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_6;
  reg [31:0] regs_7; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_7;
  reg [31:0] regs_8; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_8;
  reg [31:0] regs_9; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_9;
  reg [31:0] regs_10; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_10;
  reg [31:0] regs_11; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_11;
  reg [31:0] regs_12; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_12;
  reg [31:0] regs_13; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_13;
  reg [31:0] regs_14; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_14;
  reg [31:0] regs_15; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_15;
  reg [31:0] regs_16; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_16;
  reg [31:0] regs_17; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_17;
  reg [31:0] regs_18; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_18;
  reg [31:0] regs_19; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_19;
  reg [31:0] regs_20; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_20;
  reg [31:0] regs_21; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_21;
  reg [31:0] regs_22; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_22;
  reg [31:0] regs_23; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_23;
  reg [31:0] regs_24; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_24;
  reg [31:0] regs_25; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_25;
  reg [31:0] regs_26; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_26;
  reg [31:0] regs_27; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_27;
  reg [31:0] regs_28; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_28;
  reg [31:0] regs_29; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_29;
  reg [31:0] regs_30; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_30;
  reg [31:0] regs_31; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_31;
  reg [31:0] regs_32; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_32;
  reg [31:0] regs_33; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_33;
  reg [31:0] regs_34; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_34;
  reg [31:0] regs_35; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_35;
  reg [31:0] regs_36; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_36;
  reg [31:0] regs_37; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_37;
  reg [31:0] regs_38; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_38;
  reg [31:0] regs_39; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_39;
  reg [31:0] regs_40; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_40;
  reg [31:0] regs_41; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_41;
  reg [31:0] regs_42; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_42;
  reg [31:0] regs_43; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_43;
  reg [31:0] regs_44; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_44;
  reg [31:0] regs_45; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_45;
  reg [31:0] regs_46; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_46;
  reg [31:0] regs_47; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_47;
  reg [31:0] regs_48; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_48;
  reg [31:0] regs_49; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_49;
  reg [31:0] regs_50; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_50;
  reg [31:0] regs_51; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_51;
  reg [31:0] regs_52; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_52;
  reg [31:0] regs_53; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_53;
  reg [31:0] regs_54; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_54;
  reg [31:0] regs_55; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_55;
  reg [31:0] regs_56; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_56;
  reg [31:0] regs_57; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_57;
  reg [31:0] regs_58; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_58;
  reg [31:0] regs_59; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_59;
  reg [31:0] regs_60; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_60;
  reg [31:0] regs_61; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_61;
  reg [31:0] regs_62; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_62;
  reg [31:0] regs_63; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_63;
  reg [31:0] regs_64; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_64;
  reg [31:0] regs_65; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_65;
  reg [31:0] regs_66; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_66;
  reg [31:0] regs_67; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_67;
  reg [31:0] regs_68; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_68;
  reg [31:0] regs_69; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_69;
  reg [31:0] regs_70; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_70;
  reg [31:0] regs_71; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_71;
  reg [31:0] regs_72; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_72;
  reg [31:0] regs_73; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_73;
  reg [31:0] regs_74; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_74;
  reg [31:0] regs_75; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_75;
  reg [31:0] regs_76; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_76;
  reg [31:0] regs_77; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_77;
  reg [31:0] regs_78; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_78;
  reg [31:0] regs_79; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_79;
  reg [31:0] regs_80; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_80;
  reg [31:0] regs_81; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_81;
  reg [31:0] regs_82; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_82;
  reg [31:0] regs_83; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_83;
  reg [31:0] regs_84; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_84;
  reg [31:0] regs_85; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_85;
  reg [31:0] regs_86; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_86;
  reg [31:0] regs_87; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_87;
  reg [31:0] regs_88; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_88;
  reg [31:0] regs_89; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_89;
  reg [31:0] regs_90; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_90;
  reg [31:0] regs_91; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_91;
  reg [31:0] regs_92; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_92;
  reg [31:0] regs_93; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_93;
  reg [31:0] regs_94; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_94;
  reg [31:0] regs_95; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_95;
  reg [31:0] regs_96; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_96;
  reg [31:0] regs_97; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_97;
  reg [31:0] regs_98; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_98;
  reg [31:0] regs_99; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_99;
  assign io_out_bits_0_0 = regs_0; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_1 = regs_1; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_2 = regs_2; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_3 = regs_3; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_4 = regs_4; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_5 = regs_5; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_6 = regs_6; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_7 = regs_7; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_8 = regs_8; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_9 = regs_9; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_10 = regs_10; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_11 = regs_11; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_12 = regs_12; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_13 = regs_13; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_14 = regs_14; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_15 = regs_15; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_16 = regs_16; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_17 = regs_17; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_18 = regs_18; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_19 = regs_19; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_20 = regs_20; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_21 = regs_21; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_22 = regs_22; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_23 = regs_23; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_24 = regs_24; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_25 = regs_25; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_26 = regs_26; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_27 = regs_27; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_28 = regs_28; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_29 = regs_29; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_30 = regs_30; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_31 = regs_31; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_32 = regs_32; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_33 = regs_33; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_34 = regs_34; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_35 = regs_35; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_36 = regs_36; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_37 = regs_37; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_38 = regs_38; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_39 = regs_39; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_40 = regs_40; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_41 = regs_41; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_42 = regs_42; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_43 = regs_43; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_44 = regs_44; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_45 = regs_45; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_46 = regs_46; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_47 = regs_47; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_48 = regs_48; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_49 = regs_49; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_50 = regs_50; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_51 = regs_51; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_52 = regs_52; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_53 = regs_53; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_54 = regs_54; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_55 = regs_55; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_56 = regs_56; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_57 = regs_57; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_58 = regs_58; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_59 = regs_59; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_60 = regs_60; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_61 = regs_61; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_62 = regs_62; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_63 = regs_63; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_64 = regs_64; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_65 = regs_65; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_66 = regs_66; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_67 = regs_67; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_68 = regs_68; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_69 = regs_69; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_70 = regs_70; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_71 = regs_71; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_72 = regs_72; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_73 = regs_73; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_74 = regs_74; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_75 = regs_75; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_76 = regs_76; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_77 = regs_77; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_78 = regs_78; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_79 = regs_79; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_80 = regs_80; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_81 = regs_81; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_82 = regs_82; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_83 = regs_83; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_84 = regs_84; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_85 = regs_85; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_86 = regs_86; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_87 = regs_87; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_88 = regs_88; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_89 = regs_89; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_90 = regs_90; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_91 = regs_91; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_92 = regs_92; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_93 = regs_93; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_94 = regs_94; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_95 = regs_95; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_96 = regs_96; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_97 = regs_97; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_98 = regs_98; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_99 = regs_99; // @[MemoryBuffer.scala 65:25]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  regs_3 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  regs_4 = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  regs_5 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  regs_6 = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  regs_7 = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  regs_8 = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  regs_9 = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  regs_10 = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  regs_11 = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  regs_12 = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  regs_13 = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  regs_14 = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  regs_15 = _RAND_15[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  regs_16 = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  regs_17 = _RAND_17[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  regs_18 = _RAND_18[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  regs_19 = _RAND_19[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  regs_20 = _RAND_20[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  regs_21 = _RAND_21[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  regs_22 = _RAND_22[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  regs_23 = _RAND_23[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  regs_24 = _RAND_24[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  regs_25 = _RAND_25[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  regs_26 = _RAND_26[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  regs_27 = _RAND_27[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  regs_28 = _RAND_28[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  regs_29 = _RAND_29[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  regs_30 = _RAND_30[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  regs_31 = _RAND_31[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  regs_32 = _RAND_32[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  regs_33 = _RAND_33[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  regs_34 = _RAND_34[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  regs_35 = _RAND_35[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  regs_36 = _RAND_36[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  regs_37 = _RAND_37[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  regs_38 = _RAND_38[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  regs_39 = _RAND_39[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  regs_40 = _RAND_40[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  regs_41 = _RAND_41[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  regs_42 = _RAND_42[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  regs_43 = _RAND_43[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  regs_44 = _RAND_44[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  regs_45 = _RAND_45[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  regs_46 = _RAND_46[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  regs_47 = _RAND_47[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  regs_48 = _RAND_48[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  regs_49 = _RAND_49[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  regs_50 = _RAND_50[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  regs_51 = _RAND_51[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  regs_52 = _RAND_52[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  regs_53 = _RAND_53[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  regs_54 = _RAND_54[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  regs_55 = _RAND_55[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  regs_56 = _RAND_56[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  regs_57 = _RAND_57[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  regs_58 = _RAND_58[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  regs_59 = _RAND_59[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  regs_60 = _RAND_60[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  regs_61 = _RAND_61[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  regs_62 = _RAND_62[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  regs_63 = _RAND_63[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  regs_64 = _RAND_64[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  regs_65 = _RAND_65[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  regs_66 = _RAND_66[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  regs_67 = _RAND_67[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  regs_68 = _RAND_68[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  regs_69 = _RAND_69[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  regs_70 = _RAND_70[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  regs_71 = _RAND_71[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  regs_72 = _RAND_72[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  regs_73 = _RAND_73[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  regs_74 = _RAND_74[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  regs_75 = _RAND_75[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  regs_76 = _RAND_76[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  regs_77 = _RAND_77[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  regs_78 = _RAND_78[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  regs_79 = _RAND_79[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  regs_80 = _RAND_80[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  regs_81 = _RAND_81[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  regs_82 = _RAND_82[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  regs_83 = _RAND_83[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  regs_84 = _RAND_84[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  regs_85 = _RAND_85[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  regs_86 = _RAND_86[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  regs_87 = _RAND_87[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  regs_88 = _RAND_88[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  regs_89 = _RAND_89[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  regs_90 = _RAND_90[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  regs_91 = _RAND_91[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  regs_92 = _RAND_92[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  regs_93 = _RAND_93[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  regs_94 = _RAND_94[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  regs_95 = _RAND_95[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  regs_96 = _RAND_96[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  regs_97 = _RAND_97[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  regs_98 = _RAND_98[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  regs_99 = _RAND_99[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      regs_0 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_0 <= io_in_bits;
      end
    end
    if (reset) begin
      regs_1 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_1 <= regs_0;
      end
    end
    if (reset) begin
      regs_2 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_2 <= regs_1;
      end
    end
    if (reset) begin
      regs_3 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_3 <= regs_2;
      end
    end
    if (reset) begin
      regs_4 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_4 <= regs_3;
      end
    end
    if (reset) begin
      regs_5 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_5 <= regs_4;
      end
    end
    if (reset) begin
      regs_6 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_6 <= regs_5;
      end
    end
    if (reset) begin
      regs_7 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_7 <= regs_6;
      end
    end
    if (reset) begin
      regs_8 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_8 <= regs_7;
      end
    end
    if (reset) begin
      regs_9 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_9 <= regs_8;
      end
    end
    if (reset) begin
      regs_10 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_10 <= regs_9;
      end
    end
    if (reset) begin
      regs_11 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_11 <= regs_10;
      end
    end
    if (reset) begin
      regs_12 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_12 <= regs_11;
      end
    end
    if (reset) begin
      regs_13 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_13 <= regs_12;
      end
    end
    if (reset) begin
      regs_14 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_14 <= regs_13;
      end
    end
    if (reset) begin
      regs_15 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_15 <= regs_14;
      end
    end
    if (reset) begin
      regs_16 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_16 <= regs_15;
      end
    end
    if (reset) begin
      regs_17 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_17 <= regs_16;
      end
    end
    if (reset) begin
      regs_18 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_18 <= regs_17;
      end
    end
    if (reset) begin
      regs_19 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_19 <= regs_18;
      end
    end
    if (reset) begin
      regs_20 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_20 <= regs_19;
      end
    end
    if (reset) begin
      regs_21 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_21 <= regs_20;
      end
    end
    if (reset) begin
      regs_22 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_22 <= regs_21;
      end
    end
    if (reset) begin
      regs_23 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_23 <= regs_22;
      end
    end
    if (reset) begin
      regs_24 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_24 <= regs_23;
      end
    end
    if (reset) begin
      regs_25 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_25 <= regs_24;
      end
    end
    if (reset) begin
      regs_26 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_26 <= regs_25;
      end
    end
    if (reset) begin
      regs_27 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_27 <= regs_26;
      end
    end
    if (reset) begin
      regs_28 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_28 <= regs_27;
      end
    end
    if (reset) begin
      regs_29 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_29 <= regs_28;
      end
    end
    if (reset) begin
      regs_30 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_30 <= regs_29;
      end
    end
    if (reset) begin
      regs_31 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_31 <= regs_30;
      end
    end
    if (reset) begin
      regs_32 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_32 <= regs_31;
      end
    end
    if (reset) begin
      regs_33 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_33 <= regs_32;
      end
    end
    if (reset) begin
      regs_34 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_34 <= regs_33;
      end
    end
    if (reset) begin
      regs_35 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_35 <= regs_34;
      end
    end
    if (reset) begin
      regs_36 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_36 <= regs_35;
      end
    end
    if (reset) begin
      regs_37 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_37 <= regs_36;
      end
    end
    if (reset) begin
      regs_38 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_38 <= regs_37;
      end
    end
    if (reset) begin
      regs_39 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_39 <= regs_38;
      end
    end
    if (reset) begin
      regs_40 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_40 <= regs_39;
      end
    end
    if (reset) begin
      regs_41 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_41 <= regs_40;
      end
    end
    if (reset) begin
      regs_42 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_42 <= regs_41;
      end
    end
    if (reset) begin
      regs_43 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_43 <= regs_42;
      end
    end
    if (reset) begin
      regs_44 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_44 <= regs_43;
      end
    end
    if (reset) begin
      regs_45 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_45 <= regs_44;
      end
    end
    if (reset) begin
      regs_46 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_46 <= regs_45;
      end
    end
    if (reset) begin
      regs_47 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_47 <= regs_46;
      end
    end
    if (reset) begin
      regs_48 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_48 <= regs_47;
      end
    end
    if (reset) begin
      regs_49 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_49 <= regs_48;
      end
    end
    if (reset) begin
      regs_50 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_50 <= regs_49;
      end
    end
    if (reset) begin
      regs_51 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_51 <= regs_50;
      end
    end
    if (reset) begin
      regs_52 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_52 <= regs_51;
      end
    end
    if (reset) begin
      regs_53 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_53 <= regs_52;
      end
    end
    if (reset) begin
      regs_54 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_54 <= regs_53;
      end
    end
    if (reset) begin
      regs_55 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_55 <= regs_54;
      end
    end
    if (reset) begin
      regs_56 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_56 <= regs_55;
      end
    end
    if (reset) begin
      regs_57 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_57 <= regs_56;
      end
    end
    if (reset) begin
      regs_58 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_58 <= regs_57;
      end
    end
    if (reset) begin
      regs_59 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_59 <= regs_58;
      end
    end
    if (reset) begin
      regs_60 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_60 <= regs_59;
      end
    end
    if (reset) begin
      regs_61 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_61 <= regs_60;
      end
    end
    if (reset) begin
      regs_62 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_62 <= regs_61;
      end
    end
    if (reset) begin
      regs_63 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_63 <= regs_62;
      end
    end
    if (reset) begin
      regs_64 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_64 <= regs_63;
      end
    end
    if (reset) begin
      regs_65 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_65 <= regs_64;
      end
    end
    if (reset) begin
      regs_66 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_66 <= regs_65;
      end
    end
    if (reset) begin
      regs_67 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_67 <= regs_66;
      end
    end
    if (reset) begin
      regs_68 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_68 <= regs_67;
      end
    end
    if (reset) begin
      regs_69 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_69 <= regs_68;
      end
    end
    if (reset) begin
      regs_70 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_70 <= regs_69;
      end
    end
    if (reset) begin
      regs_71 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_71 <= regs_70;
      end
    end
    if (reset) begin
      regs_72 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_72 <= regs_71;
      end
    end
    if (reset) begin
      regs_73 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_73 <= regs_72;
      end
    end
    if (reset) begin
      regs_74 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_74 <= regs_73;
      end
    end
    if (reset) begin
      regs_75 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_75 <= regs_74;
      end
    end
    if (reset) begin
      regs_76 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_76 <= regs_75;
      end
    end
    if (reset) begin
      regs_77 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_77 <= regs_76;
      end
    end
    if (reset) begin
      regs_78 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_78 <= regs_77;
      end
    end
    if (reset) begin
      regs_79 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_79 <= regs_78;
      end
    end
    if (reset) begin
      regs_80 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_80 <= regs_79;
      end
    end
    if (reset) begin
      regs_81 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_81 <= regs_80;
      end
    end
    if (reset) begin
      regs_82 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_82 <= regs_81;
      end
    end
    if (reset) begin
      regs_83 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_83 <= regs_82;
      end
    end
    if (reset) begin
      regs_84 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_84 <= regs_83;
      end
    end
    if (reset) begin
      regs_85 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_85 <= regs_84;
      end
    end
    if (reset) begin
      regs_86 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_86 <= regs_85;
      end
    end
    if (reset) begin
      regs_87 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_87 <= regs_86;
      end
    end
    if (reset) begin
      regs_88 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_88 <= regs_87;
      end
    end
    if (reset) begin
      regs_89 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_89 <= regs_88;
      end
    end
    if (reset) begin
      regs_90 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_90 <= regs_89;
      end
    end
    if (reset) begin
      regs_91 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_91 <= regs_90;
      end
    end
    if (reset) begin
      regs_92 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_92 <= regs_91;
      end
    end
    if (reset) begin
      regs_93 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_93 <= regs_92;
      end
    end
    if (reset) begin
      regs_94 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_94 <= regs_93;
      end
    end
    if (reset) begin
      regs_95 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_95 <= regs_94;
      end
    end
    if (reset) begin
      regs_96 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_96 <= regs_95;
      end
    end
    if (reset) begin
      regs_97 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_97 <= regs_96;
      end
    end
    if (reset) begin
      regs_98 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_98 <= regs_97;
      end
    end
    if (reset) begin
      regs_99 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_99 <= regs_98;
      end
    end
  end
endmodule
module MemoryBuffer_3(
  input         clock,
  input         reset,
  input         io_in_valid,
  input  [31:0] io_in_bits,
  output [31:0] io_out_bits_0_0
);
  reg [31:0] regs_0; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_0;
  assign io_out_bits_0_0 = regs_0; // @[MemoryBuffer.scala 65:25]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      regs_0 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_0 <= io_in_bits;
      end
    end
  end
endmodule
module ConfigurationMemory(
  input         clock,
  input         reset,
  input         io_in_valid,
  input  [31:0] io_in_bits_wrdata,
  input  [2:0]  io_in_bits_wraddr,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_0_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_0_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_0_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_0_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_1_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_1_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_1_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_1_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_2_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_2_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_2_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_2_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_3_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_3_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_3_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_3_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_4_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_4_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_4_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_4_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_5_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_5_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_5_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_5_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_6_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_6_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_6_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_6_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_7_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_7_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_7_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_7_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_8_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_8_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_8_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_8_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_9_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_9_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_9_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_9_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_10_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_10_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_10_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_10_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_11_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_11_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_11_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_11_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_12_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_12_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_12_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_12_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_13_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_13_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_13_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_13_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_14_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_14_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_14_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_14_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_15_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_15_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_15_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_15_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_16_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_16_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_16_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_16_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_17_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_17_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_17_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_17_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_18_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_18_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_18_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_18_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_19_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_19_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_19_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_19_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_20_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_20_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_20_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_20_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_21_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_21_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_21_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_21_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_22_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_22_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_22_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_22_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_23_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_23_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_23_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_23_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_24_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_24_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_24_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_24_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_25_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_25_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_25_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_25_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_26_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_26_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_26_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_26_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_27_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_27_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_27_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_27_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_28_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_28_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_28_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_28_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_29_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_29_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_29_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_29_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_30_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_30_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_30_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_30_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_31_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_31_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_31_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_31_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_32_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_32_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_32_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_32_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_33_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_33_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_33_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_33_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_34_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_34_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_34_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_34_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_35_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_35_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_35_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_35_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_36_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_36_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_36_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_36_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_37_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_37_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_37_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_37_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_38_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_38_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_38_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_38_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_39_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_39_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_39_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_39_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_40_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_40_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_40_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_40_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_41_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_41_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_41_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_41_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_42_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_42_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_42_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_42_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_43_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_43_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_43_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_43_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_44_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_44_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_44_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_44_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_45_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_45_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_45_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_45_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_46_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_46_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_46_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_46_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_47_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_47_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_47_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_47_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_48_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_48_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_48_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_48_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_49_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_49_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_49_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_49_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_50_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_50_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_50_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_50_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_51_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_51_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_51_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_51_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_52_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_52_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_52_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_52_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_53_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_53_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_53_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_53_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_54_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_54_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_54_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_54_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_55_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_55_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_55_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_55_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_56_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_56_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_56_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_56_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_57_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_57_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_57_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_57_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_58_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_58_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_58_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_58_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_59_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_59_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_59_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_59_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_60_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_60_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_60_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_60_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_61_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_61_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_61_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_61_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_62_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_62_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_62_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_62_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_63_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_63_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_63_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_63_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_64_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_64_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_64_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_64_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_65_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_65_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_65_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_65_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_66_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_66_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_66_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_66_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_67_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_67_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_67_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_67_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_68_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_68_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_68_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_68_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_69_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_69_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_69_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_69_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_70_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_70_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_70_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_70_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_71_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_71_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_71_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_71_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_72_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_72_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_72_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_72_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_73_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_73_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_73_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_73_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_74_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_74_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_74_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_74_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_75_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_75_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_75_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_75_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_76_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_76_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_76_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_76_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_77_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_77_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_77_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_77_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_78_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_78_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_78_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_78_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_79_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_79_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_79_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_79_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_80_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_80_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_80_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_80_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_81_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_81_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_81_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_81_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_82_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_82_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_82_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_82_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_83_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_83_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_83_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_83_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_84_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_84_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_84_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_84_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_85_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_85_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_85_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_85_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_86_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_86_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_86_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_86_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_87_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_87_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_87_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_87_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_88_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_88_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_88_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_88_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_89_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_89_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_89_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_89_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_90_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_90_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_90_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_90_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_91_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_91_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_91_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_91_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_92_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_92_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_92_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_92_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_93_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_93_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_93_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_93_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_94_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_94_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_94_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_94_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_95_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_95_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_95_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_95_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_96_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_96_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_96_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_96_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_97_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_97_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_97_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_97_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_98_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_98_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_98_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_98_3,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_99_0,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_99_1,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_99_2,
  output [31:0] io_out_bits_confneuralNetsweightMatrix_99_3,
  output [31:0] io_out_bits_confneuralNetsweightVec_0,
  output [31:0] io_out_bits_confneuralNetsweightVec_1,
  output [31:0] io_out_bits_confneuralNetsweightVec_2,
  output [31:0] io_out_bits_confneuralNetsweightVec_3,
  output [31:0] io_out_bits_confneuralNetsweightVec_4,
  output [31:0] io_out_bits_confneuralNetsweightVec_5,
  output [31:0] io_out_bits_confneuralNetsweightVec_6,
  output [31:0] io_out_bits_confneuralNetsweightVec_7,
  output [31:0] io_out_bits_confneuralNetsweightVec_8,
  output [31:0] io_out_bits_confneuralNetsweightVec_9,
  output [31:0] io_out_bits_confneuralNetsweightVec_10,
  output [31:0] io_out_bits_confneuralNetsweightVec_11,
  output [31:0] io_out_bits_confneuralNetsweightVec_12,
  output [31:0] io_out_bits_confneuralNetsweightVec_13,
  output [31:0] io_out_bits_confneuralNetsweightVec_14,
  output [31:0] io_out_bits_confneuralNetsweightVec_15,
  output [31:0] io_out_bits_confneuralNetsweightVec_16,
  output [31:0] io_out_bits_confneuralNetsweightVec_17,
  output [31:0] io_out_bits_confneuralNetsweightVec_18,
  output [31:0] io_out_bits_confneuralNetsweightVec_19,
  output [31:0] io_out_bits_confneuralNetsweightVec_20,
  output [31:0] io_out_bits_confneuralNetsweightVec_21,
  output [31:0] io_out_bits_confneuralNetsweightVec_22,
  output [31:0] io_out_bits_confneuralNetsweightVec_23,
  output [31:0] io_out_bits_confneuralNetsweightVec_24,
  output [31:0] io_out_bits_confneuralNetsweightVec_25,
  output [31:0] io_out_bits_confneuralNetsweightVec_26,
  output [31:0] io_out_bits_confneuralNetsweightVec_27,
  output [31:0] io_out_bits_confneuralNetsweightVec_28,
  output [31:0] io_out_bits_confneuralNetsweightVec_29,
  output [31:0] io_out_bits_confneuralNetsweightVec_30,
  output [31:0] io_out_bits_confneuralNetsweightVec_31,
  output [31:0] io_out_bits_confneuralNetsweightVec_32,
  output [31:0] io_out_bits_confneuralNetsweightVec_33,
  output [31:0] io_out_bits_confneuralNetsweightVec_34,
  output [31:0] io_out_bits_confneuralNetsweightVec_35,
  output [31:0] io_out_bits_confneuralNetsweightVec_36,
  output [31:0] io_out_bits_confneuralNetsweightVec_37,
  output [31:0] io_out_bits_confneuralNetsweightVec_38,
  output [31:0] io_out_bits_confneuralNetsweightVec_39,
  output [31:0] io_out_bits_confneuralNetsweightVec_40,
  output [31:0] io_out_bits_confneuralNetsweightVec_41,
  output [31:0] io_out_bits_confneuralNetsweightVec_42,
  output [31:0] io_out_bits_confneuralNetsweightVec_43,
  output [31:0] io_out_bits_confneuralNetsweightVec_44,
  output [31:0] io_out_bits_confneuralNetsweightVec_45,
  output [31:0] io_out_bits_confneuralNetsweightVec_46,
  output [31:0] io_out_bits_confneuralNetsweightVec_47,
  output [31:0] io_out_bits_confneuralNetsweightVec_48,
  output [31:0] io_out_bits_confneuralNetsweightVec_49,
  output [31:0] io_out_bits_confneuralNetsweightVec_50,
  output [31:0] io_out_bits_confneuralNetsweightVec_51,
  output [31:0] io_out_bits_confneuralNetsweightVec_52,
  output [31:0] io_out_bits_confneuralNetsweightVec_53,
  output [31:0] io_out_bits_confneuralNetsweightVec_54,
  output [31:0] io_out_bits_confneuralNetsweightVec_55,
  output [31:0] io_out_bits_confneuralNetsweightVec_56,
  output [31:0] io_out_bits_confneuralNetsweightVec_57,
  output [31:0] io_out_bits_confneuralNetsweightVec_58,
  output [31:0] io_out_bits_confneuralNetsweightVec_59,
  output [31:0] io_out_bits_confneuralNetsweightVec_60,
  output [31:0] io_out_bits_confneuralNetsweightVec_61,
  output [31:0] io_out_bits_confneuralNetsweightVec_62,
  output [31:0] io_out_bits_confneuralNetsweightVec_63,
  output [31:0] io_out_bits_confneuralNetsweightVec_64,
  output [31:0] io_out_bits_confneuralNetsweightVec_65,
  output [31:0] io_out_bits_confneuralNetsweightVec_66,
  output [31:0] io_out_bits_confneuralNetsweightVec_67,
  output [31:0] io_out_bits_confneuralNetsweightVec_68,
  output [31:0] io_out_bits_confneuralNetsweightVec_69,
  output [31:0] io_out_bits_confneuralNetsweightVec_70,
  output [31:0] io_out_bits_confneuralNetsweightVec_71,
  output [31:0] io_out_bits_confneuralNetsweightVec_72,
  output [31:0] io_out_bits_confneuralNetsweightVec_73,
  output [31:0] io_out_bits_confneuralNetsweightVec_74,
  output [31:0] io_out_bits_confneuralNetsweightVec_75,
  output [31:0] io_out_bits_confneuralNetsweightVec_76,
  output [31:0] io_out_bits_confneuralNetsweightVec_77,
  output [31:0] io_out_bits_confneuralNetsweightVec_78,
  output [31:0] io_out_bits_confneuralNetsweightVec_79,
  output [31:0] io_out_bits_confneuralNetsweightVec_80,
  output [31:0] io_out_bits_confneuralNetsweightVec_81,
  output [31:0] io_out_bits_confneuralNetsweightVec_82,
  output [31:0] io_out_bits_confneuralNetsweightVec_83,
  output [31:0] io_out_bits_confneuralNetsweightVec_84,
  output [31:0] io_out_bits_confneuralNetsweightVec_85,
  output [31:0] io_out_bits_confneuralNetsweightVec_86,
  output [31:0] io_out_bits_confneuralNetsweightVec_87,
  output [31:0] io_out_bits_confneuralNetsweightVec_88,
  output [31:0] io_out_bits_confneuralNetsweightVec_89,
  output [31:0] io_out_bits_confneuralNetsweightVec_90,
  output [31:0] io_out_bits_confneuralNetsweightVec_91,
  output [31:0] io_out_bits_confneuralNetsweightVec_92,
  output [31:0] io_out_bits_confneuralNetsweightVec_93,
  output [31:0] io_out_bits_confneuralNetsweightVec_94,
  output [31:0] io_out_bits_confneuralNetsweightVec_95,
  output [31:0] io_out_bits_confneuralNetsweightVec_96,
  output [31:0] io_out_bits_confneuralNetsweightVec_97,
  output [31:0] io_out_bits_confneuralNetsweightVec_98,
  output [31:0] io_out_bits_confneuralNetsweightVec_99,
  output [31:0] io_out_bits_confneuralNetsbiasVec_0,
  output [31:0] io_out_bits_confneuralNetsbiasVec_1,
  output [31:0] io_out_bits_confneuralNetsbiasVec_2,
  output [31:0] io_out_bits_confneuralNetsbiasVec_3,
  output [31:0] io_out_bits_confneuralNetsbiasVec_4,
  output [31:0] io_out_bits_confneuralNetsbiasVec_5,
  output [31:0] io_out_bits_confneuralNetsbiasVec_6,
  output [31:0] io_out_bits_confneuralNetsbiasVec_7,
  output [31:0] io_out_bits_confneuralNetsbiasVec_8,
  output [31:0] io_out_bits_confneuralNetsbiasVec_9,
  output [31:0] io_out_bits_confneuralNetsbiasVec_10,
  output [31:0] io_out_bits_confneuralNetsbiasVec_11,
  output [31:0] io_out_bits_confneuralNetsbiasVec_12,
  output [31:0] io_out_bits_confneuralNetsbiasVec_13,
  output [31:0] io_out_bits_confneuralNetsbiasVec_14,
  output [31:0] io_out_bits_confneuralNetsbiasVec_15,
  output [31:0] io_out_bits_confneuralNetsbiasVec_16,
  output [31:0] io_out_bits_confneuralNetsbiasVec_17,
  output [31:0] io_out_bits_confneuralNetsbiasVec_18,
  output [31:0] io_out_bits_confneuralNetsbiasVec_19,
  output [31:0] io_out_bits_confneuralNetsbiasVec_20,
  output [31:0] io_out_bits_confneuralNetsbiasVec_21,
  output [31:0] io_out_bits_confneuralNetsbiasVec_22,
  output [31:0] io_out_bits_confneuralNetsbiasVec_23,
  output [31:0] io_out_bits_confneuralNetsbiasVec_24,
  output [31:0] io_out_bits_confneuralNetsbiasVec_25,
  output [31:0] io_out_bits_confneuralNetsbiasVec_26,
  output [31:0] io_out_bits_confneuralNetsbiasVec_27,
  output [31:0] io_out_bits_confneuralNetsbiasVec_28,
  output [31:0] io_out_bits_confneuralNetsbiasVec_29,
  output [31:0] io_out_bits_confneuralNetsbiasVec_30,
  output [31:0] io_out_bits_confneuralNetsbiasVec_31,
  output [31:0] io_out_bits_confneuralNetsbiasVec_32,
  output [31:0] io_out_bits_confneuralNetsbiasVec_33,
  output [31:0] io_out_bits_confneuralNetsbiasVec_34,
  output [31:0] io_out_bits_confneuralNetsbiasVec_35,
  output [31:0] io_out_bits_confneuralNetsbiasVec_36,
  output [31:0] io_out_bits_confneuralNetsbiasVec_37,
  output [31:0] io_out_bits_confneuralNetsbiasVec_38,
  output [31:0] io_out_bits_confneuralNetsbiasVec_39,
  output [31:0] io_out_bits_confneuralNetsbiasVec_40,
  output [31:0] io_out_bits_confneuralNetsbiasVec_41,
  output [31:0] io_out_bits_confneuralNetsbiasVec_42,
  output [31:0] io_out_bits_confneuralNetsbiasVec_43,
  output [31:0] io_out_bits_confneuralNetsbiasVec_44,
  output [31:0] io_out_bits_confneuralNetsbiasVec_45,
  output [31:0] io_out_bits_confneuralNetsbiasVec_46,
  output [31:0] io_out_bits_confneuralNetsbiasVec_47,
  output [31:0] io_out_bits_confneuralNetsbiasVec_48,
  output [31:0] io_out_bits_confneuralNetsbiasVec_49,
  output [31:0] io_out_bits_confneuralNetsbiasVec_50,
  output [31:0] io_out_bits_confneuralNetsbiasVec_51,
  output [31:0] io_out_bits_confneuralNetsbiasVec_52,
  output [31:0] io_out_bits_confneuralNetsbiasVec_53,
  output [31:0] io_out_bits_confneuralNetsbiasVec_54,
  output [31:0] io_out_bits_confneuralNetsbiasVec_55,
  output [31:0] io_out_bits_confneuralNetsbiasVec_56,
  output [31:0] io_out_bits_confneuralNetsbiasVec_57,
  output [31:0] io_out_bits_confneuralNetsbiasVec_58,
  output [31:0] io_out_bits_confneuralNetsbiasVec_59,
  output [31:0] io_out_bits_confneuralNetsbiasVec_60,
  output [31:0] io_out_bits_confneuralNetsbiasVec_61,
  output [31:0] io_out_bits_confneuralNetsbiasVec_62,
  output [31:0] io_out_bits_confneuralNetsbiasVec_63,
  output [31:0] io_out_bits_confneuralNetsbiasVec_64,
  output [31:0] io_out_bits_confneuralNetsbiasVec_65,
  output [31:0] io_out_bits_confneuralNetsbiasVec_66,
  output [31:0] io_out_bits_confneuralNetsbiasVec_67,
  output [31:0] io_out_bits_confneuralNetsbiasVec_68,
  output [31:0] io_out_bits_confneuralNetsbiasVec_69,
  output [31:0] io_out_bits_confneuralNetsbiasVec_70,
  output [31:0] io_out_bits_confneuralNetsbiasVec_71,
  output [31:0] io_out_bits_confneuralNetsbiasVec_72,
  output [31:0] io_out_bits_confneuralNetsbiasVec_73,
  output [31:0] io_out_bits_confneuralNetsbiasVec_74,
  output [31:0] io_out_bits_confneuralNetsbiasVec_75,
  output [31:0] io_out_bits_confneuralNetsbiasVec_76,
  output [31:0] io_out_bits_confneuralNetsbiasVec_77,
  output [31:0] io_out_bits_confneuralNetsbiasVec_78,
  output [31:0] io_out_bits_confneuralNetsbiasVec_79,
  output [31:0] io_out_bits_confneuralNetsbiasVec_80,
  output [31:0] io_out_bits_confneuralNetsbiasVec_81,
  output [31:0] io_out_bits_confneuralNetsbiasVec_82,
  output [31:0] io_out_bits_confneuralNetsbiasVec_83,
  output [31:0] io_out_bits_confneuralNetsbiasVec_84,
  output [31:0] io_out_bits_confneuralNetsbiasVec_85,
  output [31:0] io_out_bits_confneuralNetsbiasVec_86,
  output [31:0] io_out_bits_confneuralNetsbiasVec_87,
  output [31:0] io_out_bits_confneuralNetsbiasVec_88,
  output [31:0] io_out_bits_confneuralNetsbiasVec_89,
  output [31:0] io_out_bits_confneuralNetsbiasVec_90,
  output [31:0] io_out_bits_confneuralNetsbiasVec_91,
  output [31:0] io_out_bits_confneuralNetsbiasVec_92,
  output [31:0] io_out_bits_confneuralNetsbiasVec_93,
  output [31:0] io_out_bits_confneuralNetsbiasVec_94,
  output [31:0] io_out_bits_confneuralNetsbiasVec_95,
  output [31:0] io_out_bits_confneuralNetsbiasVec_96,
  output [31:0] io_out_bits_confneuralNetsbiasVec_97,
  output [31:0] io_out_bits_confneuralNetsbiasVec_98,
  output [31:0] io_out_bits_confneuralNetsbiasVec_99,
  output [31:0] io_out_bits_confneuralNetsbiasScalar_0,
  output        io_out_bits_confInputMuxSel
);
  wire  neuralNetsweightMatrixMemory_clock; // @[ConfigurationMemory.scala 60:44]
  wire  neuralNetsweightMatrixMemory_reset; // @[ConfigurationMemory.scala 60:44]
  wire  neuralNetsweightMatrixMemory_io_in_valid; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_in_bits; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_0_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_0_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_0_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_0_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_1_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_1_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_1_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_1_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_2_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_2_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_2_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_2_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_3_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_3_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_3_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_3_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_4_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_4_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_4_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_4_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_5_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_5_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_5_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_5_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_6_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_6_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_6_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_6_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_7_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_7_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_7_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_7_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_8_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_8_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_8_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_8_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_9_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_9_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_9_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_9_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_10_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_10_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_10_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_10_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_11_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_11_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_11_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_11_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_12_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_12_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_12_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_12_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_13_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_13_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_13_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_13_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_14_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_14_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_14_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_14_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_15_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_15_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_15_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_15_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_16_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_16_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_16_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_16_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_17_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_17_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_17_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_17_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_18_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_18_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_18_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_18_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_19_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_19_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_19_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_19_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_20_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_20_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_20_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_20_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_21_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_21_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_21_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_21_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_22_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_22_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_22_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_22_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_23_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_23_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_23_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_23_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_24_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_24_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_24_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_24_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_25_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_25_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_25_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_25_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_26_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_26_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_26_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_26_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_27_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_27_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_27_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_27_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_28_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_28_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_28_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_28_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_29_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_29_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_29_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_29_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_30_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_30_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_30_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_30_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_31_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_31_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_31_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_31_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_32_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_32_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_32_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_32_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_33_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_33_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_33_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_33_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_34_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_34_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_34_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_34_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_35_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_35_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_35_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_35_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_36_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_36_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_36_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_36_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_37_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_37_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_37_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_37_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_38_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_38_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_38_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_38_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_39_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_39_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_39_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_39_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_40_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_40_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_40_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_40_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_41_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_41_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_41_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_41_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_42_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_42_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_42_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_42_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_43_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_43_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_43_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_43_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_44_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_44_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_44_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_44_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_45_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_45_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_45_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_45_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_46_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_46_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_46_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_46_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_47_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_47_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_47_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_47_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_48_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_48_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_48_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_48_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_49_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_49_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_49_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_49_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_50_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_50_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_50_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_50_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_51_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_51_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_51_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_51_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_52_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_52_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_52_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_52_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_53_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_53_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_53_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_53_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_54_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_54_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_54_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_54_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_55_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_55_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_55_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_55_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_56_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_56_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_56_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_56_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_57_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_57_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_57_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_57_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_58_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_58_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_58_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_58_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_59_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_59_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_59_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_59_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_60_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_60_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_60_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_60_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_61_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_61_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_61_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_61_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_62_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_62_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_62_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_62_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_63_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_63_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_63_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_63_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_64_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_64_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_64_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_64_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_65_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_65_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_65_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_65_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_66_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_66_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_66_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_66_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_67_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_67_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_67_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_67_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_68_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_68_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_68_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_68_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_69_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_69_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_69_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_69_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_70_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_70_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_70_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_70_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_71_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_71_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_71_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_71_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_72_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_72_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_72_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_72_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_73_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_73_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_73_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_73_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_74_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_74_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_74_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_74_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_75_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_75_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_75_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_75_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_76_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_76_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_76_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_76_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_77_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_77_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_77_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_77_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_78_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_78_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_78_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_78_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_79_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_79_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_79_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_79_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_80_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_80_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_80_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_80_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_81_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_81_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_81_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_81_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_82_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_82_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_82_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_82_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_83_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_83_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_83_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_83_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_84_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_84_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_84_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_84_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_85_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_85_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_85_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_85_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_86_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_86_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_86_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_86_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_87_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_87_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_87_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_87_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_88_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_88_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_88_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_88_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_89_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_89_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_89_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_89_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_90_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_90_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_90_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_90_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_91_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_91_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_91_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_91_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_92_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_92_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_92_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_92_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_93_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_93_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_93_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_93_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_94_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_94_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_94_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_94_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_95_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_95_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_95_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_95_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_96_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_96_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_96_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_96_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_97_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_97_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_97_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_97_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_98_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_98_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_98_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_98_3; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_99_0; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_99_1; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_99_2; // @[ConfigurationMemory.scala 60:44]
  wire [31:0] neuralNetsweightMatrixMemory_io_out_bits_99_3; // @[ConfigurationMemory.scala 60:44]
  wire  neuralNetsweightVecMemory_clock; // @[ConfigurationMemory.scala 72:41]
  wire  neuralNetsweightVecMemory_reset; // @[ConfigurationMemory.scala 72:41]
  wire  neuralNetsweightVecMemory_io_in_valid; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_in_bits; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_0; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_1; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_2; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_3; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_4; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_5; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_6; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_7; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_8; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_9; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_10; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_11; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_12; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_13; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_14; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_15; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_16; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_17; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_18; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_19; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_20; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_21; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_22; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_23; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_24; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_25; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_26; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_27; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_28; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_29; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_30; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_31; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_32; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_33; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_34; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_35; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_36; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_37; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_38; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_39; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_40; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_41; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_42; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_43; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_44; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_45; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_46; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_47; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_48; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_49; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_50; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_51; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_52; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_53; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_54; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_55; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_56; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_57; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_58; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_59; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_60; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_61; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_62; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_63; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_64; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_65; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_66; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_67; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_68; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_69; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_70; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_71; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_72; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_73; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_74; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_75; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_76; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_77; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_78; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_79; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_80; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_81; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_82; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_83; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_84; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_85; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_86; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_87; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_88; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_89; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_90; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_91; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_92; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_93; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_94; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_95; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_96; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_97; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_98; // @[ConfigurationMemory.scala 72:41]
  wire [31:0] neuralNetsweightVecMemory_io_out_bits_0_99; // @[ConfigurationMemory.scala 72:41]
  wire  neuralNetsbiasVecMemory_clock; // @[ConfigurationMemory.scala 83:39]
  wire  neuralNetsbiasVecMemory_reset; // @[ConfigurationMemory.scala 83:39]
  wire  neuralNetsbiasVecMemory_io_in_valid; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_in_bits; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_0; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_1; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_2; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_3; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_4; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_5; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_6; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_7; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_8; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_9; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_10; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_11; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_12; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_13; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_14; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_15; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_16; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_17; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_18; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_19; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_20; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_21; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_22; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_23; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_24; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_25; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_26; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_27; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_28; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_29; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_30; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_31; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_32; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_33; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_34; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_35; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_36; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_37; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_38; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_39; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_40; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_41; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_42; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_43; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_44; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_45; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_46; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_47; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_48; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_49; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_50; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_51; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_52; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_53; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_54; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_55; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_56; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_57; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_58; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_59; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_60; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_61; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_62; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_63; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_64; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_65; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_66; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_67; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_68; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_69; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_70; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_71; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_72; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_73; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_74; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_75; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_76; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_77; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_78; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_79; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_80; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_81; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_82; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_83; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_84; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_85; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_86; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_87; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_88; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_89; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_90; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_91; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_92; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_93; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_94; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_95; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_96; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_97; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_98; // @[ConfigurationMemory.scala 83:39]
  wire [31:0] neuralNetsbiasVecMemory_io_out_bits_0_99; // @[ConfigurationMemory.scala 83:39]
  wire  neuralNetsbiasScalarMemory_clock; // @[ConfigurationMemory.scala 95:42]
  wire  neuralNetsbiasScalarMemory_reset; // @[ConfigurationMemory.scala 95:42]
  wire  neuralNetsbiasScalarMemory_io_in_valid; // @[ConfigurationMemory.scala 95:42]
  wire [31:0] neuralNetsbiasScalarMemory_io_in_bits; // @[ConfigurationMemory.scala 95:42]
  wire [31:0] neuralNetsbiasScalarMemory_io_out_bits_0_0; // @[ConfigurationMemory.scala 95:42]
  wire  _T; // @[ConfigurationMemory.scala 63:68]
  wire  _T_2; // @[ConfigurationMemory.scala 75:65]
  wire  _T_4; // @[ConfigurationMemory.scala 86:63]
  wire  _T_6; // @[ConfigurationMemory.scala 98:66]
  reg  inputMuxSel; // @[ConfigurationMemory.scala 103:28]
  reg [31:0] _RAND_0;
  wire  _T_8; // @[ConfigurationMemory.scala 104:29]
  wire  _T_9; // @[ConfigurationMemory.scala 104:20]
  wire [31:0] _T_10; // @[ConfigurationMemory.scala 104:90]
  wire  _T_11; // @[ConfigurationMemory.scala 104:92]
  MemoryBuffer neuralNetsweightMatrixMemory ( // @[ConfigurationMemory.scala 60:44]
    .clock(neuralNetsweightMatrixMemory_clock),
    .reset(neuralNetsweightMatrixMemory_reset),
    .io_in_valid(neuralNetsweightMatrixMemory_io_in_valid),
    .io_in_bits(neuralNetsweightMatrixMemory_io_in_bits),
    .io_out_bits_0_0(neuralNetsweightMatrixMemory_io_out_bits_0_0),
    .io_out_bits_0_1(neuralNetsweightMatrixMemory_io_out_bits_0_1),
    .io_out_bits_0_2(neuralNetsweightMatrixMemory_io_out_bits_0_2),
    .io_out_bits_0_3(neuralNetsweightMatrixMemory_io_out_bits_0_3),
    .io_out_bits_1_0(neuralNetsweightMatrixMemory_io_out_bits_1_0),
    .io_out_bits_1_1(neuralNetsweightMatrixMemory_io_out_bits_1_1),
    .io_out_bits_1_2(neuralNetsweightMatrixMemory_io_out_bits_1_2),
    .io_out_bits_1_3(neuralNetsweightMatrixMemory_io_out_bits_1_3),
    .io_out_bits_2_0(neuralNetsweightMatrixMemory_io_out_bits_2_0),
    .io_out_bits_2_1(neuralNetsweightMatrixMemory_io_out_bits_2_1),
    .io_out_bits_2_2(neuralNetsweightMatrixMemory_io_out_bits_2_2),
    .io_out_bits_2_3(neuralNetsweightMatrixMemory_io_out_bits_2_3),
    .io_out_bits_3_0(neuralNetsweightMatrixMemory_io_out_bits_3_0),
    .io_out_bits_3_1(neuralNetsweightMatrixMemory_io_out_bits_3_1),
    .io_out_bits_3_2(neuralNetsweightMatrixMemory_io_out_bits_3_2),
    .io_out_bits_3_3(neuralNetsweightMatrixMemory_io_out_bits_3_3),
    .io_out_bits_4_0(neuralNetsweightMatrixMemory_io_out_bits_4_0),
    .io_out_bits_4_1(neuralNetsweightMatrixMemory_io_out_bits_4_1),
    .io_out_bits_4_2(neuralNetsweightMatrixMemory_io_out_bits_4_2),
    .io_out_bits_4_3(neuralNetsweightMatrixMemory_io_out_bits_4_3),
    .io_out_bits_5_0(neuralNetsweightMatrixMemory_io_out_bits_5_0),
    .io_out_bits_5_1(neuralNetsweightMatrixMemory_io_out_bits_5_1),
    .io_out_bits_5_2(neuralNetsweightMatrixMemory_io_out_bits_5_2),
    .io_out_bits_5_3(neuralNetsweightMatrixMemory_io_out_bits_5_3),
    .io_out_bits_6_0(neuralNetsweightMatrixMemory_io_out_bits_6_0),
    .io_out_bits_6_1(neuralNetsweightMatrixMemory_io_out_bits_6_1),
    .io_out_bits_6_2(neuralNetsweightMatrixMemory_io_out_bits_6_2),
    .io_out_bits_6_3(neuralNetsweightMatrixMemory_io_out_bits_6_3),
    .io_out_bits_7_0(neuralNetsweightMatrixMemory_io_out_bits_7_0),
    .io_out_bits_7_1(neuralNetsweightMatrixMemory_io_out_bits_7_1),
    .io_out_bits_7_2(neuralNetsweightMatrixMemory_io_out_bits_7_2),
    .io_out_bits_7_3(neuralNetsweightMatrixMemory_io_out_bits_7_3),
    .io_out_bits_8_0(neuralNetsweightMatrixMemory_io_out_bits_8_0),
    .io_out_bits_8_1(neuralNetsweightMatrixMemory_io_out_bits_8_1),
    .io_out_bits_8_2(neuralNetsweightMatrixMemory_io_out_bits_8_2),
    .io_out_bits_8_3(neuralNetsweightMatrixMemory_io_out_bits_8_3),
    .io_out_bits_9_0(neuralNetsweightMatrixMemory_io_out_bits_9_0),
    .io_out_bits_9_1(neuralNetsweightMatrixMemory_io_out_bits_9_1),
    .io_out_bits_9_2(neuralNetsweightMatrixMemory_io_out_bits_9_2),
    .io_out_bits_9_3(neuralNetsweightMatrixMemory_io_out_bits_9_3),
    .io_out_bits_10_0(neuralNetsweightMatrixMemory_io_out_bits_10_0),
    .io_out_bits_10_1(neuralNetsweightMatrixMemory_io_out_bits_10_1),
    .io_out_bits_10_2(neuralNetsweightMatrixMemory_io_out_bits_10_2),
    .io_out_bits_10_3(neuralNetsweightMatrixMemory_io_out_bits_10_3),
    .io_out_bits_11_0(neuralNetsweightMatrixMemory_io_out_bits_11_0),
    .io_out_bits_11_1(neuralNetsweightMatrixMemory_io_out_bits_11_1),
    .io_out_bits_11_2(neuralNetsweightMatrixMemory_io_out_bits_11_2),
    .io_out_bits_11_3(neuralNetsweightMatrixMemory_io_out_bits_11_3),
    .io_out_bits_12_0(neuralNetsweightMatrixMemory_io_out_bits_12_0),
    .io_out_bits_12_1(neuralNetsweightMatrixMemory_io_out_bits_12_1),
    .io_out_bits_12_2(neuralNetsweightMatrixMemory_io_out_bits_12_2),
    .io_out_bits_12_3(neuralNetsweightMatrixMemory_io_out_bits_12_3),
    .io_out_bits_13_0(neuralNetsweightMatrixMemory_io_out_bits_13_0),
    .io_out_bits_13_1(neuralNetsweightMatrixMemory_io_out_bits_13_1),
    .io_out_bits_13_2(neuralNetsweightMatrixMemory_io_out_bits_13_2),
    .io_out_bits_13_3(neuralNetsweightMatrixMemory_io_out_bits_13_3),
    .io_out_bits_14_0(neuralNetsweightMatrixMemory_io_out_bits_14_0),
    .io_out_bits_14_1(neuralNetsweightMatrixMemory_io_out_bits_14_1),
    .io_out_bits_14_2(neuralNetsweightMatrixMemory_io_out_bits_14_2),
    .io_out_bits_14_3(neuralNetsweightMatrixMemory_io_out_bits_14_3),
    .io_out_bits_15_0(neuralNetsweightMatrixMemory_io_out_bits_15_0),
    .io_out_bits_15_1(neuralNetsweightMatrixMemory_io_out_bits_15_1),
    .io_out_bits_15_2(neuralNetsweightMatrixMemory_io_out_bits_15_2),
    .io_out_bits_15_3(neuralNetsweightMatrixMemory_io_out_bits_15_3),
    .io_out_bits_16_0(neuralNetsweightMatrixMemory_io_out_bits_16_0),
    .io_out_bits_16_1(neuralNetsweightMatrixMemory_io_out_bits_16_1),
    .io_out_bits_16_2(neuralNetsweightMatrixMemory_io_out_bits_16_2),
    .io_out_bits_16_3(neuralNetsweightMatrixMemory_io_out_bits_16_3),
    .io_out_bits_17_0(neuralNetsweightMatrixMemory_io_out_bits_17_0),
    .io_out_bits_17_1(neuralNetsweightMatrixMemory_io_out_bits_17_1),
    .io_out_bits_17_2(neuralNetsweightMatrixMemory_io_out_bits_17_2),
    .io_out_bits_17_3(neuralNetsweightMatrixMemory_io_out_bits_17_3),
    .io_out_bits_18_0(neuralNetsweightMatrixMemory_io_out_bits_18_0),
    .io_out_bits_18_1(neuralNetsweightMatrixMemory_io_out_bits_18_1),
    .io_out_bits_18_2(neuralNetsweightMatrixMemory_io_out_bits_18_2),
    .io_out_bits_18_3(neuralNetsweightMatrixMemory_io_out_bits_18_3),
    .io_out_bits_19_0(neuralNetsweightMatrixMemory_io_out_bits_19_0),
    .io_out_bits_19_1(neuralNetsweightMatrixMemory_io_out_bits_19_1),
    .io_out_bits_19_2(neuralNetsweightMatrixMemory_io_out_bits_19_2),
    .io_out_bits_19_3(neuralNetsweightMatrixMemory_io_out_bits_19_3),
    .io_out_bits_20_0(neuralNetsweightMatrixMemory_io_out_bits_20_0),
    .io_out_bits_20_1(neuralNetsweightMatrixMemory_io_out_bits_20_1),
    .io_out_bits_20_2(neuralNetsweightMatrixMemory_io_out_bits_20_2),
    .io_out_bits_20_3(neuralNetsweightMatrixMemory_io_out_bits_20_3),
    .io_out_bits_21_0(neuralNetsweightMatrixMemory_io_out_bits_21_0),
    .io_out_bits_21_1(neuralNetsweightMatrixMemory_io_out_bits_21_1),
    .io_out_bits_21_2(neuralNetsweightMatrixMemory_io_out_bits_21_2),
    .io_out_bits_21_3(neuralNetsweightMatrixMemory_io_out_bits_21_3),
    .io_out_bits_22_0(neuralNetsweightMatrixMemory_io_out_bits_22_0),
    .io_out_bits_22_1(neuralNetsweightMatrixMemory_io_out_bits_22_1),
    .io_out_bits_22_2(neuralNetsweightMatrixMemory_io_out_bits_22_2),
    .io_out_bits_22_3(neuralNetsweightMatrixMemory_io_out_bits_22_3),
    .io_out_bits_23_0(neuralNetsweightMatrixMemory_io_out_bits_23_0),
    .io_out_bits_23_1(neuralNetsweightMatrixMemory_io_out_bits_23_1),
    .io_out_bits_23_2(neuralNetsweightMatrixMemory_io_out_bits_23_2),
    .io_out_bits_23_3(neuralNetsweightMatrixMemory_io_out_bits_23_3),
    .io_out_bits_24_0(neuralNetsweightMatrixMemory_io_out_bits_24_0),
    .io_out_bits_24_1(neuralNetsweightMatrixMemory_io_out_bits_24_1),
    .io_out_bits_24_2(neuralNetsweightMatrixMemory_io_out_bits_24_2),
    .io_out_bits_24_3(neuralNetsweightMatrixMemory_io_out_bits_24_3),
    .io_out_bits_25_0(neuralNetsweightMatrixMemory_io_out_bits_25_0),
    .io_out_bits_25_1(neuralNetsweightMatrixMemory_io_out_bits_25_1),
    .io_out_bits_25_2(neuralNetsweightMatrixMemory_io_out_bits_25_2),
    .io_out_bits_25_3(neuralNetsweightMatrixMemory_io_out_bits_25_3),
    .io_out_bits_26_0(neuralNetsweightMatrixMemory_io_out_bits_26_0),
    .io_out_bits_26_1(neuralNetsweightMatrixMemory_io_out_bits_26_1),
    .io_out_bits_26_2(neuralNetsweightMatrixMemory_io_out_bits_26_2),
    .io_out_bits_26_3(neuralNetsweightMatrixMemory_io_out_bits_26_3),
    .io_out_bits_27_0(neuralNetsweightMatrixMemory_io_out_bits_27_0),
    .io_out_bits_27_1(neuralNetsweightMatrixMemory_io_out_bits_27_1),
    .io_out_bits_27_2(neuralNetsweightMatrixMemory_io_out_bits_27_2),
    .io_out_bits_27_3(neuralNetsweightMatrixMemory_io_out_bits_27_3),
    .io_out_bits_28_0(neuralNetsweightMatrixMemory_io_out_bits_28_0),
    .io_out_bits_28_1(neuralNetsweightMatrixMemory_io_out_bits_28_1),
    .io_out_bits_28_2(neuralNetsweightMatrixMemory_io_out_bits_28_2),
    .io_out_bits_28_3(neuralNetsweightMatrixMemory_io_out_bits_28_3),
    .io_out_bits_29_0(neuralNetsweightMatrixMemory_io_out_bits_29_0),
    .io_out_bits_29_1(neuralNetsweightMatrixMemory_io_out_bits_29_1),
    .io_out_bits_29_2(neuralNetsweightMatrixMemory_io_out_bits_29_2),
    .io_out_bits_29_3(neuralNetsweightMatrixMemory_io_out_bits_29_3),
    .io_out_bits_30_0(neuralNetsweightMatrixMemory_io_out_bits_30_0),
    .io_out_bits_30_1(neuralNetsweightMatrixMemory_io_out_bits_30_1),
    .io_out_bits_30_2(neuralNetsweightMatrixMemory_io_out_bits_30_2),
    .io_out_bits_30_3(neuralNetsweightMatrixMemory_io_out_bits_30_3),
    .io_out_bits_31_0(neuralNetsweightMatrixMemory_io_out_bits_31_0),
    .io_out_bits_31_1(neuralNetsweightMatrixMemory_io_out_bits_31_1),
    .io_out_bits_31_2(neuralNetsweightMatrixMemory_io_out_bits_31_2),
    .io_out_bits_31_3(neuralNetsweightMatrixMemory_io_out_bits_31_3),
    .io_out_bits_32_0(neuralNetsweightMatrixMemory_io_out_bits_32_0),
    .io_out_bits_32_1(neuralNetsweightMatrixMemory_io_out_bits_32_1),
    .io_out_bits_32_2(neuralNetsweightMatrixMemory_io_out_bits_32_2),
    .io_out_bits_32_3(neuralNetsweightMatrixMemory_io_out_bits_32_3),
    .io_out_bits_33_0(neuralNetsweightMatrixMemory_io_out_bits_33_0),
    .io_out_bits_33_1(neuralNetsweightMatrixMemory_io_out_bits_33_1),
    .io_out_bits_33_2(neuralNetsweightMatrixMemory_io_out_bits_33_2),
    .io_out_bits_33_3(neuralNetsweightMatrixMemory_io_out_bits_33_3),
    .io_out_bits_34_0(neuralNetsweightMatrixMemory_io_out_bits_34_0),
    .io_out_bits_34_1(neuralNetsweightMatrixMemory_io_out_bits_34_1),
    .io_out_bits_34_2(neuralNetsweightMatrixMemory_io_out_bits_34_2),
    .io_out_bits_34_3(neuralNetsweightMatrixMemory_io_out_bits_34_3),
    .io_out_bits_35_0(neuralNetsweightMatrixMemory_io_out_bits_35_0),
    .io_out_bits_35_1(neuralNetsweightMatrixMemory_io_out_bits_35_1),
    .io_out_bits_35_2(neuralNetsweightMatrixMemory_io_out_bits_35_2),
    .io_out_bits_35_3(neuralNetsweightMatrixMemory_io_out_bits_35_3),
    .io_out_bits_36_0(neuralNetsweightMatrixMemory_io_out_bits_36_0),
    .io_out_bits_36_1(neuralNetsweightMatrixMemory_io_out_bits_36_1),
    .io_out_bits_36_2(neuralNetsweightMatrixMemory_io_out_bits_36_2),
    .io_out_bits_36_3(neuralNetsweightMatrixMemory_io_out_bits_36_3),
    .io_out_bits_37_0(neuralNetsweightMatrixMemory_io_out_bits_37_0),
    .io_out_bits_37_1(neuralNetsweightMatrixMemory_io_out_bits_37_1),
    .io_out_bits_37_2(neuralNetsweightMatrixMemory_io_out_bits_37_2),
    .io_out_bits_37_3(neuralNetsweightMatrixMemory_io_out_bits_37_3),
    .io_out_bits_38_0(neuralNetsweightMatrixMemory_io_out_bits_38_0),
    .io_out_bits_38_1(neuralNetsweightMatrixMemory_io_out_bits_38_1),
    .io_out_bits_38_2(neuralNetsweightMatrixMemory_io_out_bits_38_2),
    .io_out_bits_38_3(neuralNetsweightMatrixMemory_io_out_bits_38_3),
    .io_out_bits_39_0(neuralNetsweightMatrixMemory_io_out_bits_39_0),
    .io_out_bits_39_1(neuralNetsweightMatrixMemory_io_out_bits_39_1),
    .io_out_bits_39_2(neuralNetsweightMatrixMemory_io_out_bits_39_2),
    .io_out_bits_39_3(neuralNetsweightMatrixMemory_io_out_bits_39_3),
    .io_out_bits_40_0(neuralNetsweightMatrixMemory_io_out_bits_40_0),
    .io_out_bits_40_1(neuralNetsweightMatrixMemory_io_out_bits_40_1),
    .io_out_bits_40_2(neuralNetsweightMatrixMemory_io_out_bits_40_2),
    .io_out_bits_40_3(neuralNetsweightMatrixMemory_io_out_bits_40_3),
    .io_out_bits_41_0(neuralNetsweightMatrixMemory_io_out_bits_41_0),
    .io_out_bits_41_1(neuralNetsweightMatrixMemory_io_out_bits_41_1),
    .io_out_bits_41_2(neuralNetsweightMatrixMemory_io_out_bits_41_2),
    .io_out_bits_41_3(neuralNetsweightMatrixMemory_io_out_bits_41_3),
    .io_out_bits_42_0(neuralNetsweightMatrixMemory_io_out_bits_42_0),
    .io_out_bits_42_1(neuralNetsweightMatrixMemory_io_out_bits_42_1),
    .io_out_bits_42_2(neuralNetsweightMatrixMemory_io_out_bits_42_2),
    .io_out_bits_42_3(neuralNetsweightMatrixMemory_io_out_bits_42_3),
    .io_out_bits_43_0(neuralNetsweightMatrixMemory_io_out_bits_43_0),
    .io_out_bits_43_1(neuralNetsweightMatrixMemory_io_out_bits_43_1),
    .io_out_bits_43_2(neuralNetsweightMatrixMemory_io_out_bits_43_2),
    .io_out_bits_43_3(neuralNetsweightMatrixMemory_io_out_bits_43_3),
    .io_out_bits_44_0(neuralNetsweightMatrixMemory_io_out_bits_44_0),
    .io_out_bits_44_1(neuralNetsweightMatrixMemory_io_out_bits_44_1),
    .io_out_bits_44_2(neuralNetsweightMatrixMemory_io_out_bits_44_2),
    .io_out_bits_44_3(neuralNetsweightMatrixMemory_io_out_bits_44_3),
    .io_out_bits_45_0(neuralNetsweightMatrixMemory_io_out_bits_45_0),
    .io_out_bits_45_1(neuralNetsweightMatrixMemory_io_out_bits_45_1),
    .io_out_bits_45_2(neuralNetsweightMatrixMemory_io_out_bits_45_2),
    .io_out_bits_45_3(neuralNetsweightMatrixMemory_io_out_bits_45_3),
    .io_out_bits_46_0(neuralNetsweightMatrixMemory_io_out_bits_46_0),
    .io_out_bits_46_1(neuralNetsweightMatrixMemory_io_out_bits_46_1),
    .io_out_bits_46_2(neuralNetsweightMatrixMemory_io_out_bits_46_2),
    .io_out_bits_46_3(neuralNetsweightMatrixMemory_io_out_bits_46_3),
    .io_out_bits_47_0(neuralNetsweightMatrixMemory_io_out_bits_47_0),
    .io_out_bits_47_1(neuralNetsweightMatrixMemory_io_out_bits_47_1),
    .io_out_bits_47_2(neuralNetsweightMatrixMemory_io_out_bits_47_2),
    .io_out_bits_47_3(neuralNetsweightMatrixMemory_io_out_bits_47_3),
    .io_out_bits_48_0(neuralNetsweightMatrixMemory_io_out_bits_48_0),
    .io_out_bits_48_1(neuralNetsweightMatrixMemory_io_out_bits_48_1),
    .io_out_bits_48_2(neuralNetsweightMatrixMemory_io_out_bits_48_2),
    .io_out_bits_48_3(neuralNetsweightMatrixMemory_io_out_bits_48_3),
    .io_out_bits_49_0(neuralNetsweightMatrixMemory_io_out_bits_49_0),
    .io_out_bits_49_1(neuralNetsweightMatrixMemory_io_out_bits_49_1),
    .io_out_bits_49_2(neuralNetsweightMatrixMemory_io_out_bits_49_2),
    .io_out_bits_49_3(neuralNetsweightMatrixMemory_io_out_bits_49_3),
    .io_out_bits_50_0(neuralNetsweightMatrixMemory_io_out_bits_50_0),
    .io_out_bits_50_1(neuralNetsweightMatrixMemory_io_out_bits_50_1),
    .io_out_bits_50_2(neuralNetsweightMatrixMemory_io_out_bits_50_2),
    .io_out_bits_50_3(neuralNetsweightMatrixMemory_io_out_bits_50_3),
    .io_out_bits_51_0(neuralNetsweightMatrixMemory_io_out_bits_51_0),
    .io_out_bits_51_1(neuralNetsweightMatrixMemory_io_out_bits_51_1),
    .io_out_bits_51_2(neuralNetsweightMatrixMemory_io_out_bits_51_2),
    .io_out_bits_51_3(neuralNetsweightMatrixMemory_io_out_bits_51_3),
    .io_out_bits_52_0(neuralNetsweightMatrixMemory_io_out_bits_52_0),
    .io_out_bits_52_1(neuralNetsweightMatrixMemory_io_out_bits_52_1),
    .io_out_bits_52_2(neuralNetsweightMatrixMemory_io_out_bits_52_2),
    .io_out_bits_52_3(neuralNetsweightMatrixMemory_io_out_bits_52_3),
    .io_out_bits_53_0(neuralNetsweightMatrixMemory_io_out_bits_53_0),
    .io_out_bits_53_1(neuralNetsweightMatrixMemory_io_out_bits_53_1),
    .io_out_bits_53_2(neuralNetsweightMatrixMemory_io_out_bits_53_2),
    .io_out_bits_53_3(neuralNetsweightMatrixMemory_io_out_bits_53_3),
    .io_out_bits_54_0(neuralNetsweightMatrixMemory_io_out_bits_54_0),
    .io_out_bits_54_1(neuralNetsweightMatrixMemory_io_out_bits_54_1),
    .io_out_bits_54_2(neuralNetsweightMatrixMemory_io_out_bits_54_2),
    .io_out_bits_54_3(neuralNetsweightMatrixMemory_io_out_bits_54_3),
    .io_out_bits_55_0(neuralNetsweightMatrixMemory_io_out_bits_55_0),
    .io_out_bits_55_1(neuralNetsweightMatrixMemory_io_out_bits_55_1),
    .io_out_bits_55_2(neuralNetsweightMatrixMemory_io_out_bits_55_2),
    .io_out_bits_55_3(neuralNetsweightMatrixMemory_io_out_bits_55_3),
    .io_out_bits_56_0(neuralNetsweightMatrixMemory_io_out_bits_56_0),
    .io_out_bits_56_1(neuralNetsweightMatrixMemory_io_out_bits_56_1),
    .io_out_bits_56_2(neuralNetsweightMatrixMemory_io_out_bits_56_2),
    .io_out_bits_56_3(neuralNetsweightMatrixMemory_io_out_bits_56_3),
    .io_out_bits_57_0(neuralNetsweightMatrixMemory_io_out_bits_57_0),
    .io_out_bits_57_1(neuralNetsweightMatrixMemory_io_out_bits_57_1),
    .io_out_bits_57_2(neuralNetsweightMatrixMemory_io_out_bits_57_2),
    .io_out_bits_57_3(neuralNetsweightMatrixMemory_io_out_bits_57_3),
    .io_out_bits_58_0(neuralNetsweightMatrixMemory_io_out_bits_58_0),
    .io_out_bits_58_1(neuralNetsweightMatrixMemory_io_out_bits_58_1),
    .io_out_bits_58_2(neuralNetsweightMatrixMemory_io_out_bits_58_2),
    .io_out_bits_58_3(neuralNetsweightMatrixMemory_io_out_bits_58_3),
    .io_out_bits_59_0(neuralNetsweightMatrixMemory_io_out_bits_59_0),
    .io_out_bits_59_1(neuralNetsweightMatrixMemory_io_out_bits_59_1),
    .io_out_bits_59_2(neuralNetsweightMatrixMemory_io_out_bits_59_2),
    .io_out_bits_59_3(neuralNetsweightMatrixMemory_io_out_bits_59_3),
    .io_out_bits_60_0(neuralNetsweightMatrixMemory_io_out_bits_60_0),
    .io_out_bits_60_1(neuralNetsweightMatrixMemory_io_out_bits_60_1),
    .io_out_bits_60_2(neuralNetsweightMatrixMemory_io_out_bits_60_2),
    .io_out_bits_60_3(neuralNetsweightMatrixMemory_io_out_bits_60_3),
    .io_out_bits_61_0(neuralNetsweightMatrixMemory_io_out_bits_61_0),
    .io_out_bits_61_1(neuralNetsweightMatrixMemory_io_out_bits_61_1),
    .io_out_bits_61_2(neuralNetsweightMatrixMemory_io_out_bits_61_2),
    .io_out_bits_61_3(neuralNetsweightMatrixMemory_io_out_bits_61_3),
    .io_out_bits_62_0(neuralNetsweightMatrixMemory_io_out_bits_62_0),
    .io_out_bits_62_1(neuralNetsweightMatrixMemory_io_out_bits_62_1),
    .io_out_bits_62_2(neuralNetsweightMatrixMemory_io_out_bits_62_2),
    .io_out_bits_62_3(neuralNetsweightMatrixMemory_io_out_bits_62_3),
    .io_out_bits_63_0(neuralNetsweightMatrixMemory_io_out_bits_63_0),
    .io_out_bits_63_1(neuralNetsweightMatrixMemory_io_out_bits_63_1),
    .io_out_bits_63_2(neuralNetsweightMatrixMemory_io_out_bits_63_2),
    .io_out_bits_63_3(neuralNetsweightMatrixMemory_io_out_bits_63_3),
    .io_out_bits_64_0(neuralNetsweightMatrixMemory_io_out_bits_64_0),
    .io_out_bits_64_1(neuralNetsweightMatrixMemory_io_out_bits_64_1),
    .io_out_bits_64_2(neuralNetsweightMatrixMemory_io_out_bits_64_2),
    .io_out_bits_64_3(neuralNetsweightMatrixMemory_io_out_bits_64_3),
    .io_out_bits_65_0(neuralNetsweightMatrixMemory_io_out_bits_65_0),
    .io_out_bits_65_1(neuralNetsweightMatrixMemory_io_out_bits_65_1),
    .io_out_bits_65_2(neuralNetsweightMatrixMemory_io_out_bits_65_2),
    .io_out_bits_65_3(neuralNetsweightMatrixMemory_io_out_bits_65_3),
    .io_out_bits_66_0(neuralNetsweightMatrixMemory_io_out_bits_66_0),
    .io_out_bits_66_1(neuralNetsweightMatrixMemory_io_out_bits_66_1),
    .io_out_bits_66_2(neuralNetsweightMatrixMemory_io_out_bits_66_2),
    .io_out_bits_66_3(neuralNetsweightMatrixMemory_io_out_bits_66_3),
    .io_out_bits_67_0(neuralNetsweightMatrixMemory_io_out_bits_67_0),
    .io_out_bits_67_1(neuralNetsweightMatrixMemory_io_out_bits_67_1),
    .io_out_bits_67_2(neuralNetsweightMatrixMemory_io_out_bits_67_2),
    .io_out_bits_67_3(neuralNetsweightMatrixMemory_io_out_bits_67_3),
    .io_out_bits_68_0(neuralNetsweightMatrixMemory_io_out_bits_68_0),
    .io_out_bits_68_1(neuralNetsweightMatrixMemory_io_out_bits_68_1),
    .io_out_bits_68_2(neuralNetsweightMatrixMemory_io_out_bits_68_2),
    .io_out_bits_68_3(neuralNetsweightMatrixMemory_io_out_bits_68_3),
    .io_out_bits_69_0(neuralNetsweightMatrixMemory_io_out_bits_69_0),
    .io_out_bits_69_1(neuralNetsweightMatrixMemory_io_out_bits_69_1),
    .io_out_bits_69_2(neuralNetsweightMatrixMemory_io_out_bits_69_2),
    .io_out_bits_69_3(neuralNetsweightMatrixMemory_io_out_bits_69_3),
    .io_out_bits_70_0(neuralNetsweightMatrixMemory_io_out_bits_70_0),
    .io_out_bits_70_1(neuralNetsweightMatrixMemory_io_out_bits_70_1),
    .io_out_bits_70_2(neuralNetsweightMatrixMemory_io_out_bits_70_2),
    .io_out_bits_70_3(neuralNetsweightMatrixMemory_io_out_bits_70_3),
    .io_out_bits_71_0(neuralNetsweightMatrixMemory_io_out_bits_71_0),
    .io_out_bits_71_1(neuralNetsweightMatrixMemory_io_out_bits_71_1),
    .io_out_bits_71_2(neuralNetsweightMatrixMemory_io_out_bits_71_2),
    .io_out_bits_71_3(neuralNetsweightMatrixMemory_io_out_bits_71_3),
    .io_out_bits_72_0(neuralNetsweightMatrixMemory_io_out_bits_72_0),
    .io_out_bits_72_1(neuralNetsweightMatrixMemory_io_out_bits_72_1),
    .io_out_bits_72_2(neuralNetsweightMatrixMemory_io_out_bits_72_2),
    .io_out_bits_72_3(neuralNetsweightMatrixMemory_io_out_bits_72_3),
    .io_out_bits_73_0(neuralNetsweightMatrixMemory_io_out_bits_73_0),
    .io_out_bits_73_1(neuralNetsweightMatrixMemory_io_out_bits_73_1),
    .io_out_bits_73_2(neuralNetsweightMatrixMemory_io_out_bits_73_2),
    .io_out_bits_73_3(neuralNetsweightMatrixMemory_io_out_bits_73_3),
    .io_out_bits_74_0(neuralNetsweightMatrixMemory_io_out_bits_74_0),
    .io_out_bits_74_1(neuralNetsweightMatrixMemory_io_out_bits_74_1),
    .io_out_bits_74_2(neuralNetsweightMatrixMemory_io_out_bits_74_2),
    .io_out_bits_74_3(neuralNetsweightMatrixMemory_io_out_bits_74_3),
    .io_out_bits_75_0(neuralNetsweightMatrixMemory_io_out_bits_75_0),
    .io_out_bits_75_1(neuralNetsweightMatrixMemory_io_out_bits_75_1),
    .io_out_bits_75_2(neuralNetsweightMatrixMemory_io_out_bits_75_2),
    .io_out_bits_75_3(neuralNetsweightMatrixMemory_io_out_bits_75_3),
    .io_out_bits_76_0(neuralNetsweightMatrixMemory_io_out_bits_76_0),
    .io_out_bits_76_1(neuralNetsweightMatrixMemory_io_out_bits_76_1),
    .io_out_bits_76_2(neuralNetsweightMatrixMemory_io_out_bits_76_2),
    .io_out_bits_76_3(neuralNetsweightMatrixMemory_io_out_bits_76_3),
    .io_out_bits_77_0(neuralNetsweightMatrixMemory_io_out_bits_77_0),
    .io_out_bits_77_1(neuralNetsweightMatrixMemory_io_out_bits_77_1),
    .io_out_bits_77_2(neuralNetsweightMatrixMemory_io_out_bits_77_2),
    .io_out_bits_77_3(neuralNetsweightMatrixMemory_io_out_bits_77_3),
    .io_out_bits_78_0(neuralNetsweightMatrixMemory_io_out_bits_78_0),
    .io_out_bits_78_1(neuralNetsweightMatrixMemory_io_out_bits_78_1),
    .io_out_bits_78_2(neuralNetsweightMatrixMemory_io_out_bits_78_2),
    .io_out_bits_78_3(neuralNetsweightMatrixMemory_io_out_bits_78_3),
    .io_out_bits_79_0(neuralNetsweightMatrixMemory_io_out_bits_79_0),
    .io_out_bits_79_1(neuralNetsweightMatrixMemory_io_out_bits_79_1),
    .io_out_bits_79_2(neuralNetsweightMatrixMemory_io_out_bits_79_2),
    .io_out_bits_79_3(neuralNetsweightMatrixMemory_io_out_bits_79_3),
    .io_out_bits_80_0(neuralNetsweightMatrixMemory_io_out_bits_80_0),
    .io_out_bits_80_1(neuralNetsweightMatrixMemory_io_out_bits_80_1),
    .io_out_bits_80_2(neuralNetsweightMatrixMemory_io_out_bits_80_2),
    .io_out_bits_80_3(neuralNetsweightMatrixMemory_io_out_bits_80_3),
    .io_out_bits_81_0(neuralNetsweightMatrixMemory_io_out_bits_81_0),
    .io_out_bits_81_1(neuralNetsweightMatrixMemory_io_out_bits_81_1),
    .io_out_bits_81_2(neuralNetsweightMatrixMemory_io_out_bits_81_2),
    .io_out_bits_81_3(neuralNetsweightMatrixMemory_io_out_bits_81_3),
    .io_out_bits_82_0(neuralNetsweightMatrixMemory_io_out_bits_82_0),
    .io_out_bits_82_1(neuralNetsweightMatrixMemory_io_out_bits_82_1),
    .io_out_bits_82_2(neuralNetsweightMatrixMemory_io_out_bits_82_2),
    .io_out_bits_82_3(neuralNetsweightMatrixMemory_io_out_bits_82_3),
    .io_out_bits_83_0(neuralNetsweightMatrixMemory_io_out_bits_83_0),
    .io_out_bits_83_1(neuralNetsweightMatrixMemory_io_out_bits_83_1),
    .io_out_bits_83_2(neuralNetsweightMatrixMemory_io_out_bits_83_2),
    .io_out_bits_83_3(neuralNetsweightMatrixMemory_io_out_bits_83_3),
    .io_out_bits_84_0(neuralNetsweightMatrixMemory_io_out_bits_84_0),
    .io_out_bits_84_1(neuralNetsweightMatrixMemory_io_out_bits_84_1),
    .io_out_bits_84_2(neuralNetsweightMatrixMemory_io_out_bits_84_2),
    .io_out_bits_84_3(neuralNetsweightMatrixMemory_io_out_bits_84_3),
    .io_out_bits_85_0(neuralNetsweightMatrixMemory_io_out_bits_85_0),
    .io_out_bits_85_1(neuralNetsweightMatrixMemory_io_out_bits_85_1),
    .io_out_bits_85_2(neuralNetsweightMatrixMemory_io_out_bits_85_2),
    .io_out_bits_85_3(neuralNetsweightMatrixMemory_io_out_bits_85_3),
    .io_out_bits_86_0(neuralNetsweightMatrixMemory_io_out_bits_86_0),
    .io_out_bits_86_1(neuralNetsweightMatrixMemory_io_out_bits_86_1),
    .io_out_bits_86_2(neuralNetsweightMatrixMemory_io_out_bits_86_2),
    .io_out_bits_86_3(neuralNetsweightMatrixMemory_io_out_bits_86_3),
    .io_out_bits_87_0(neuralNetsweightMatrixMemory_io_out_bits_87_0),
    .io_out_bits_87_1(neuralNetsweightMatrixMemory_io_out_bits_87_1),
    .io_out_bits_87_2(neuralNetsweightMatrixMemory_io_out_bits_87_2),
    .io_out_bits_87_3(neuralNetsweightMatrixMemory_io_out_bits_87_3),
    .io_out_bits_88_0(neuralNetsweightMatrixMemory_io_out_bits_88_0),
    .io_out_bits_88_1(neuralNetsweightMatrixMemory_io_out_bits_88_1),
    .io_out_bits_88_2(neuralNetsweightMatrixMemory_io_out_bits_88_2),
    .io_out_bits_88_3(neuralNetsweightMatrixMemory_io_out_bits_88_3),
    .io_out_bits_89_0(neuralNetsweightMatrixMemory_io_out_bits_89_0),
    .io_out_bits_89_1(neuralNetsweightMatrixMemory_io_out_bits_89_1),
    .io_out_bits_89_2(neuralNetsweightMatrixMemory_io_out_bits_89_2),
    .io_out_bits_89_3(neuralNetsweightMatrixMemory_io_out_bits_89_3),
    .io_out_bits_90_0(neuralNetsweightMatrixMemory_io_out_bits_90_0),
    .io_out_bits_90_1(neuralNetsweightMatrixMemory_io_out_bits_90_1),
    .io_out_bits_90_2(neuralNetsweightMatrixMemory_io_out_bits_90_2),
    .io_out_bits_90_3(neuralNetsweightMatrixMemory_io_out_bits_90_3),
    .io_out_bits_91_0(neuralNetsweightMatrixMemory_io_out_bits_91_0),
    .io_out_bits_91_1(neuralNetsweightMatrixMemory_io_out_bits_91_1),
    .io_out_bits_91_2(neuralNetsweightMatrixMemory_io_out_bits_91_2),
    .io_out_bits_91_3(neuralNetsweightMatrixMemory_io_out_bits_91_3),
    .io_out_bits_92_0(neuralNetsweightMatrixMemory_io_out_bits_92_0),
    .io_out_bits_92_1(neuralNetsweightMatrixMemory_io_out_bits_92_1),
    .io_out_bits_92_2(neuralNetsweightMatrixMemory_io_out_bits_92_2),
    .io_out_bits_92_3(neuralNetsweightMatrixMemory_io_out_bits_92_3),
    .io_out_bits_93_0(neuralNetsweightMatrixMemory_io_out_bits_93_0),
    .io_out_bits_93_1(neuralNetsweightMatrixMemory_io_out_bits_93_1),
    .io_out_bits_93_2(neuralNetsweightMatrixMemory_io_out_bits_93_2),
    .io_out_bits_93_3(neuralNetsweightMatrixMemory_io_out_bits_93_3),
    .io_out_bits_94_0(neuralNetsweightMatrixMemory_io_out_bits_94_0),
    .io_out_bits_94_1(neuralNetsweightMatrixMemory_io_out_bits_94_1),
    .io_out_bits_94_2(neuralNetsweightMatrixMemory_io_out_bits_94_2),
    .io_out_bits_94_3(neuralNetsweightMatrixMemory_io_out_bits_94_3),
    .io_out_bits_95_0(neuralNetsweightMatrixMemory_io_out_bits_95_0),
    .io_out_bits_95_1(neuralNetsweightMatrixMemory_io_out_bits_95_1),
    .io_out_bits_95_2(neuralNetsweightMatrixMemory_io_out_bits_95_2),
    .io_out_bits_95_3(neuralNetsweightMatrixMemory_io_out_bits_95_3),
    .io_out_bits_96_0(neuralNetsweightMatrixMemory_io_out_bits_96_0),
    .io_out_bits_96_1(neuralNetsweightMatrixMemory_io_out_bits_96_1),
    .io_out_bits_96_2(neuralNetsweightMatrixMemory_io_out_bits_96_2),
    .io_out_bits_96_3(neuralNetsweightMatrixMemory_io_out_bits_96_3),
    .io_out_bits_97_0(neuralNetsweightMatrixMemory_io_out_bits_97_0),
    .io_out_bits_97_1(neuralNetsweightMatrixMemory_io_out_bits_97_1),
    .io_out_bits_97_2(neuralNetsweightMatrixMemory_io_out_bits_97_2),
    .io_out_bits_97_3(neuralNetsweightMatrixMemory_io_out_bits_97_3),
    .io_out_bits_98_0(neuralNetsweightMatrixMemory_io_out_bits_98_0),
    .io_out_bits_98_1(neuralNetsweightMatrixMemory_io_out_bits_98_1),
    .io_out_bits_98_2(neuralNetsweightMatrixMemory_io_out_bits_98_2),
    .io_out_bits_98_3(neuralNetsweightMatrixMemory_io_out_bits_98_3),
    .io_out_bits_99_0(neuralNetsweightMatrixMemory_io_out_bits_99_0),
    .io_out_bits_99_1(neuralNetsweightMatrixMemory_io_out_bits_99_1),
    .io_out_bits_99_2(neuralNetsweightMatrixMemory_io_out_bits_99_2),
    .io_out_bits_99_3(neuralNetsweightMatrixMemory_io_out_bits_99_3)
  );
  MemoryBuffer_1 neuralNetsweightVecMemory ( // @[ConfigurationMemory.scala 72:41]
    .clock(neuralNetsweightVecMemory_clock),
    .reset(neuralNetsweightVecMemory_reset),
    .io_in_valid(neuralNetsweightVecMemory_io_in_valid),
    .io_in_bits(neuralNetsweightVecMemory_io_in_bits),
    .io_out_bits_0_0(neuralNetsweightVecMemory_io_out_bits_0_0),
    .io_out_bits_0_1(neuralNetsweightVecMemory_io_out_bits_0_1),
    .io_out_bits_0_2(neuralNetsweightVecMemory_io_out_bits_0_2),
    .io_out_bits_0_3(neuralNetsweightVecMemory_io_out_bits_0_3),
    .io_out_bits_0_4(neuralNetsweightVecMemory_io_out_bits_0_4),
    .io_out_bits_0_5(neuralNetsweightVecMemory_io_out_bits_0_5),
    .io_out_bits_0_6(neuralNetsweightVecMemory_io_out_bits_0_6),
    .io_out_bits_0_7(neuralNetsweightVecMemory_io_out_bits_0_7),
    .io_out_bits_0_8(neuralNetsweightVecMemory_io_out_bits_0_8),
    .io_out_bits_0_9(neuralNetsweightVecMemory_io_out_bits_0_9),
    .io_out_bits_0_10(neuralNetsweightVecMemory_io_out_bits_0_10),
    .io_out_bits_0_11(neuralNetsweightVecMemory_io_out_bits_0_11),
    .io_out_bits_0_12(neuralNetsweightVecMemory_io_out_bits_0_12),
    .io_out_bits_0_13(neuralNetsweightVecMemory_io_out_bits_0_13),
    .io_out_bits_0_14(neuralNetsweightVecMemory_io_out_bits_0_14),
    .io_out_bits_0_15(neuralNetsweightVecMemory_io_out_bits_0_15),
    .io_out_bits_0_16(neuralNetsweightVecMemory_io_out_bits_0_16),
    .io_out_bits_0_17(neuralNetsweightVecMemory_io_out_bits_0_17),
    .io_out_bits_0_18(neuralNetsweightVecMemory_io_out_bits_0_18),
    .io_out_bits_0_19(neuralNetsweightVecMemory_io_out_bits_0_19),
    .io_out_bits_0_20(neuralNetsweightVecMemory_io_out_bits_0_20),
    .io_out_bits_0_21(neuralNetsweightVecMemory_io_out_bits_0_21),
    .io_out_bits_0_22(neuralNetsweightVecMemory_io_out_bits_0_22),
    .io_out_bits_0_23(neuralNetsweightVecMemory_io_out_bits_0_23),
    .io_out_bits_0_24(neuralNetsweightVecMemory_io_out_bits_0_24),
    .io_out_bits_0_25(neuralNetsweightVecMemory_io_out_bits_0_25),
    .io_out_bits_0_26(neuralNetsweightVecMemory_io_out_bits_0_26),
    .io_out_bits_0_27(neuralNetsweightVecMemory_io_out_bits_0_27),
    .io_out_bits_0_28(neuralNetsweightVecMemory_io_out_bits_0_28),
    .io_out_bits_0_29(neuralNetsweightVecMemory_io_out_bits_0_29),
    .io_out_bits_0_30(neuralNetsweightVecMemory_io_out_bits_0_30),
    .io_out_bits_0_31(neuralNetsweightVecMemory_io_out_bits_0_31),
    .io_out_bits_0_32(neuralNetsweightVecMemory_io_out_bits_0_32),
    .io_out_bits_0_33(neuralNetsweightVecMemory_io_out_bits_0_33),
    .io_out_bits_0_34(neuralNetsweightVecMemory_io_out_bits_0_34),
    .io_out_bits_0_35(neuralNetsweightVecMemory_io_out_bits_0_35),
    .io_out_bits_0_36(neuralNetsweightVecMemory_io_out_bits_0_36),
    .io_out_bits_0_37(neuralNetsweightVecMemory_io_out_bits_0_37),
    .io_out_bits_0_38(neuralNetsweightVecMemory_io_out_bits_0_38),
    .io_out_bits_0_39(neuralNetsweightVecMemory_io_out_bits_0_39),
    .io_out_bits_0_40(neuralNetsweightVecMemory_io_out_bits_0_40),
    .io_out_bits_0_41(neuralNetsweightVecMemory_io_out_bits_0_41),
    .io_out_bits_0_42(neuralNetsweightVecMemory_io_out_bits_0_42),
    .io_out_bits_0_43(neuralNetsweightVecMemory_io_out_bits_0_43),
    .io_out_bits_0_44(neuralNetsweightVecMemory_io_out_bits_0_44),
    .io_out_bits_0_45(neuralNetsweightVecMemory_io_out_bits_0_45),
    .io_out_bits_0_46(neuralNetsweightVecMemory_io_out_bits_0_46),
    .io_out_bits_0_47(neuralNetsweightVecMemory_io_out_bits_0_47),
    .io_out_bits_0_48(neuralNetsweightVecMemory_io_out_bits_0_48),
    .io_out_bits_0_49(neuralNetsweightVecMemory_io_out_bits_0_49),
    .io_out_bits_0_50(neuralNetsweightVecMemory_io_out_bits_0_50),
    .io_out_bits_0_51(neuralNetsweightVecMemory_io_out_bits_0_51),
    .io_out_bits_0_52(neuralNetsweightVecMemory_io_out_bits_0_52),
    .io_out_bits_0_53(neuralNetsweightVecMemory_io_out_bits_0_53),
    .io_out_bits_0_54(neuralNetsweightVecMemory_io_out_bits_0_54),
    .io_out_bits_0_55(neuralNetsweightVecMemory_io_out_bits_0_55),
    .io_out_bits_0_56(neuralNetsweightVecMemory_io_out_bits_0_56),
    .io_out_bits_0_57(neuralNetsweightVecMemory_io_out_bits_0_57),
    .io_out_bits_0_58(neuralNetsweightVecMemory_io_out_bits_0_58),
    .io_out_bits_0_59(neuralNetsweightVecMemory_io_out_bits_0_59),
    .io_out_bits_0_60(neuralNetsweightVecMemory_io_out_bits_0_60),
    .io_out_bits_0_61(neuralNetsweightVecMemory_io_out_bits_0_61),
    .io_out_bits_0_62(neuralNetsweightVecMemory_io_out_bits_0_62),
    .io_out_bits_0_63(neuralNetsweightVecMemory_io_out_bits_0_63),
    .io_out_bits_0_64(neuralNetsweightVecMemory_io_out_bits_0_64),
    .io_out_bits_0_65(neuralNetsweightVecMemory_io_out_bits_0_65),
    .io_out_bits_0_66(neuralNetsweightVecMemory_io_out_bits_0_66),
    .io_out_bits_0_67(neuralNetsweightVecMemory_io_out_bits_0_67),
    .io_out_bits_0_68(neuralNetsweightVecMemory_io_out_bits_0_68),
    .io_out_bits_0_69(neuralNetsweightVecMemory_io_out_bits_0_69),
    .io_out_bits_0_70(neuralNetsweightVecMemory_io_out_bits_0_70),
    .io_out_bits_0_71(neuralNetsweightVecMemory_io_out_bits_0_71),
    .io_out_bits_0_72(neuralNetsweightVecMemory_io_out_bits_0_72),
    .io_out_bits_0_73(neuralNetsweightVecMemory_io_out_bits_0_73),
    .io_out_bits_0_74(neuralNetsweightVecMemory_io_out_bits_0_74),
    .io_out_bits_0_75(neuralNetsweightVecMemory_io_out_bits_0_75),
    .io_out_bits_0_76(neuralNetsweightVecMemory_io_out_bits_0_76),
    .io_out_bits_0_77(neuralNetsweightVecMemory_io_out_bits_0_77),
    .io_out_bits_0_78(neuralNetsweightVecMemory_io_out_bits_0_78),
    .io_out_bits_0_79(neuralNetsweightVecMemory_io_out_bits_0_79),
    .io_out_bits_0_80(neuralNetsweightVecMemory_io_out_bits_0_80),
    .io_out_bits_0_81(neuralNetsweightVecMemory_io_out_bits_0_81),
    .io_out_bits_0_82(neuralNetsweightVecMemory_io_out_bits_0_82),
    .io_out_bits_0_83(neuralNetsweightVecMemory_io_out_bits_0_83),
    .io_out_bits_0_84(neuralNetsweightVecMemory_io_out_bits_0_84),
    .io_out_bits_0_85(neuralNetsweightVecMemory_io_out_bits_0_85),
    .io_out_bits_0_86(neuralNetsweightVecMemory_io_out_bits_0_86),
    .io_out_bits_0_87(neuralNetsweightVecMemory_io_out_bits_0_87),
    .io_out_bits_0_88(neuralNetsweightVecMemory_io_out_bits_0_88),
    .io_out_bits_0_89(neuralNetsweightVecMemory_io_out_bits_0_89),
    .io_out_bits_0_90(neuralNetsweightVecMemory_io_out_bits_0_90),
    .io_out_bits_0_91(neuralNetsweightVecMemory_io_out_bits_0_91),
    .io_out_bits_0_92(neuralNetsweightVecMemory_io_out_bits_0_92),
    .io_out_bits_0_93(neuralNetsweightVecMemory_io_out_bits_0_93),
    .io_out_bits_0_94(neuralNetsweightVecMemory_io_out_bits_0_94),
    .io_out_bits_0_95(neuralNetsweightVecMemory_io_out_bits_0_95),
    .io_out_bits_0_96(neuralNetsweightVecMemory_io_out_bits_0_96),
    .io_out_bits_0_97(neuralNetsweightVecMemory_io_out_bits_0_97),
    .io_out_bits_0_98(neuralNetsweightVecMemory_io_out_bits_0_98),
    .io_out_bits_0_99(neuralNetsweightVecMemory_io_out_bits_0_99)
  );
  MemoryBuffer_1 neuralNetsbiasVecMemory ( // @[ConfigurationMemory.scala 83:39]
    .clock(neuralNetsbiasVecMemory_clock),
    .reset(neuralNetsbiasVecMemory_reset),
    .io_in_valid(neuralNetsbiasVecMemory_io_in_valid),
    .io_in_bits(neuralNetsbiasVecMemory_io_in_bits),
    .io_out_bits_0_0(neuralNetsbiasVecMemory_io_out_bits_0_0),
    .io_out_bits_0_1(neuralNetsbiasVecMemory_io_out_bits_0_1),
    .io_out_bits_0_2(neuralNetsbiasVecMemory_io_out_bits_0_2),
    .io_out_bits_0_3(neuralNetsbiasVecMemory_io_out_bits_0_3),
    .io_out_bits_0_4(neuralNetsbiasVecMemory_io_out_bits_0_4),
    .io_out_bits_0_5(neuralNetsbiasVecMemory_io_out_bits_0_5),
    .io_out_bits_0_6(neuralNetsbiasVecMemory_io_out_bits_0_6),
    .io_out_bits_0_7(neuralNetsbiasVecMemory_io_out_bits_0_7),
    .io_out_bits_0_8(neuralNetsbiasVecMemory_io_out_bits_0_8),
    .io_out_bits_0_9(neuralNetsbiasVecMemory_io_out_bits_0_9),
    .io_out_bits_0_10(neuralNetsbiasVecMemory_io_out_bits_0_10),
    .io_out_bits_0_11(neuralNetsbiasVecMemory_io_out_bits_0_11),
    .io_out_bits_0_12(neuralNetsbiasVecMemory_io_out_bits_0_12),
    .io_out_bits_0_13(neuralNetsbiasVecMemory_io_out_bits_0_13),
    .io_out_bits_0_14(neuralNetsbiasVecMemory_io_out_bits_0_14),
    .io_out_bits_0_15(neuralNetsbiasVecMemory_io_out_bits_0_15),
    .io_out_bits_0_16(neuralNetsbiasVecMemory_io_out_bits_0_16),
    .io_out_bits_0_17(neuralNetsbiasVecMemory_io_out_bits_0_17),
    .io_out_bits_0_18(neuralNetsbiasVecMemory_io_out_bits_0_18),
    .io_out_bits_0_19(neuralNetsbiasVecMemory_io_out_bits_0_19),
    .io_out_bits_0_20(neuralNetsbiasVecMemory_io_out_bits_0_20),
    .io_out_bits_0_21(neuralNetsbiasVecMemory_io_out_bits_0_21),
    .io_out_bits_0_22(neuralNetsbiasVecMemory_io_out_bits_0_22),
    .io_out_bits_0_23(neuralNetsbiasVecMemory_io_out_bits_0_23),
    .io_out_bits_0_24(neuralNetsbiasVecMemory_io_out_bits_0_24),
    .io_out_bits_0_25(neuralNetsbiasVecMemory_io_out_bits_0_25),
    .io_out_bits_0_26(neuralNetsbiasVecMemory_io_out_bits_0_26),
    .io_out_bits_0_27(neuralNetsbiasVecMemory_io_out_bits_0_27),
    .io_out_bits_0_28(neuralNetsbiasVecMemory_io_out_bits_0_28),
    .io_out_bits_0_29(neuralNetsbiasVecMemory_io_out_bits_0_29),
    .io_out_bits_0_30(neuralNetsbiasVecMemory_io_out_bits_0_30),
    .io_out_bits_0_31(neuralNetsbiasVecMemory_io_out_bits_0_31),
    .io_out_bits_0_32(neuralNetsbiasVecMemory_io_out_bits_0_32),
    .io_out_bits_0_33(neuralNetsbiasVecMemory_io_out_bits_0_33),
    .io_out_bits_0_34(neuralNetsbiasVecMemory_io_out_bits_0_34),
    .io_out_bits_0_35(neuralNetsbiasVecMemory_io_out_bits_0_35),
    .io_out_bits_0_36(neuralNetsbiasVecMemory_io_out_bits_0_36),
    .io_out_bits_0_37(neuralNetsbiasVecMemory_io_out_bits_0_37),
    .io_out_bits_0_38(neuralNetsbiasVecMemory_io_out_bits_0_38),
    .io_out_bits_0_39(neuralNetsbiasVecMemory_io_out_bits_0_39),
    .io_out_bits_0_40(neuralNetsbiasVecMemory_io_out_bits_0_40),
    .io_out_bits_0_41(neuralNetsbiasVecMemory_io_out_bits_0_41),
    .io_out_bits_0_42(neuralNetsbiasVecMemory_io_out_bits_0_42),
    .io_out_bits_0_43(neuralNetsbiasVecMemory_io_out_bits_0_43),
    .io_out_bits_0_44(neuralNetsbiasVecMemory_io_out_bits_0_44),
    .io_out_bits_0_45(neuralNetsbiasVecMemory_io_out_bits_0_45),
    .io_out_bits_0_46(neuralNetsbiasVecMemory_io_out_bits_0_46),
    .io_out_bits_0_47(neuralNetsbiasVecMemory_io_out_bits_0_47),
    .io_out_bits_0_48(neuralNetsbiasVecMemory_io_out_bits_0_48),
    .io_out_bits_0_49(neuralNetsbiasVecMemory_io_out_bits_0_49),
    .io_out_bits_0_50(neuralNetsbiasVecMemory_io_out_bits_0_50),
    .io_out_bits_0_51(neuralNetsbiasVecMemory_io_out_bits_0_51),
    .io_out_bits_0_52(neuralNetsbiasVecMemory_io_out_bits_0_52),
    .io_out_bits_0_53(neuralNetsbiasVecMemory_io_out_bits_0_53),
    .io_out_bits_0_54(neuralNetsbiasVecMemory_io_out_bits_0_54),
    .io_out_bits_0_55(neuralNetsbiasVecMemory_io_out_bits_0_55),
    .io_out_bits_0_56(neuralNetsbiasVecMemory_io_out_bits_0_56),
    .io_out_bits_0_57(neuralNetsbiasVecMemory_io_out_bits_0_57),
    .io_out_bits_0_58(neuralNetsbiasVecMemory_io_out_bits_0_58),
    .io_out_bits_0_59(neuralNetsbiasVecMemory_io_out_bits_0_59),
    .io_out_bits_0_60(neuralNetsbiasVecMemory_io_out_bits_0_60),
    .io_out_bits_0_61(neuralNetsbiasVecMemory_io_out_bits_0_61),
    .io_out_bits_0_62(neuralNetsbiasVecMemory_io_out_bits_0_62),
    .io_out_bits_0_63(neuralNetsbiasVecMemory_io_out_bits_0_63),
    .io_out_bits_0_64(neuralNetsbiasVecMemory_io_out_bits_0_64),
    .io_out_bits_0_65(neuralNetsbiasVecMemory_io_out_bits_0_65),
    .io_out_bits_0_66(neuralNetsbiasVecMemory_io_out_bits_0_66),
    .io_out_bits_0_67(neuralNetsbiasVecMemory_io_out_bits_0_67),
    .io_out_bits_0_68(neuralNetsbiasVecMemory_io_out_bits_0_68),
    .io_out_bits_0_69(neuralNetsbiasVecMemory_io_out_bits_0_69),
    .io_out_bits_0_70(neuralNetsbiasVecMemory_io_out_bits_0_70),
    .io_out_bits_0_71(neuralNetsbiasVecMemory_io_out_bits_0_71),
    .io_out_bits_0_72(neuralNetsbiasVecMemory_io_out_bits_0_72),
    .io_out_bits_0_73(neuralNetsbiasVecMemory_io_out_bits_0_73),
    .io_out_bits_0_74(neuralNetsbiasVecMemory_io_out_bits_0_74),
    .io_out_bits_0_75(neuralNetsbiasVecMemory_io_out_bits_0_75),
    .io_out_bits_0_76(neuralNetsbiasVecMemory_io_out_bits_0_76),
    .io_out_bits_0_77(neuralNetsbiasVecMemory_io_out_bits_0_77),
    .io_out_bits_0_78(neuralNetsbiasVecMemory_io_out_bits_0_78),
    .io_out_bits_0_79(neuralNetsbiasVecMemory_io_out_bits_0_79),
    .io_out_bits_0_80(neuralNetsbiasVecMemory_io_out_bits_0_80),
    .io_out_bits_0_81(neuralNetsbiasVecMemory_io_out_bits_0_81),
    .io_out_bits_0_82(neuralNetsbiasVecMemory_io_out_bits_0_82),
    .io_out_bits_0_83(neuralNetsbiasVecMemory_io_out_bits_0_83),
    .io_out_bits_0_84(neuralNetsbiasVecMemory_io_out_bits_0_84),
    .io_out_bits_0_85(neuralNetsbiasVecMemory_io_out_bits_0_85),
    .io_out_bits_0_86(neuralNetsbiasVecMemory_io_out_bits_0_86),
    .io_out_bits_0_87(neuralNetsbiasVecMemory_io_out_bits_0_87),
    .io_out_bits_0_88(neuralNetsbiasVecMemory_io_out_bits_0_88),
    .io_out_bits_0_89(neuralNetsbiasVecMemory_io_out_bits_0_89),
    .io_out_bits_0_90(neuralNetsbiasVecMemory_io_out_bits_0_90),
    .io_out_bits_0_91(neuralNetsbiasVecMemory_io_out_bits_0_91),
    .io_out_bits_0_92(neuralNetsbiasVecMemory_io_out_bits_0_92),
    .io_out_bits_0_93(neuralNetsbiasVecMemory_io_out_bits_0_93),
    .io_out_bits_0_94(neuralNetsbiasVecMemory_io_out_bits_0_94),
    .io_out_bits_0_95(neuralNetsbiasVecMemory_io_out_bits_0_95),
    .io_out_bits_0_96(neuralNetsbiasVecMemory_io_out_bits_0_96),
    .io_out_bits_0_97(neuralNetsbiasVecMemory_io_out_bits_0_97),
    .io_out_bits_0_98(neuralNetsbiasVecMemory_io_out_bits_0_98),
    .io_out_bits_0_99(neuralNetsbiasVecMemory_io_out_bits_0_99)
  );
  MemoryBuffer_3 neuralNetsbiasScalarMemory ( // @[ConfigurationMemory.scala 95:42]
    .clock(neuralNetsbiasScalarMemory_clock),
    .reset(neuralNetsbiasScalarMemory_reset),
    .io_in_valid(neuralNetsbiasScalarMemory_io_in_valid),
    .io_in_bits(neuralNetsbiasScalarMemory_io_in_bits),
    .io_out_bits_0_0(neuralNetsbiasScalarMemory_io_out_bits_0_0)
  );
  assign _T = io_in_bits_wraddr == 3'h0; // @[ConfigurationMemory.scala 63:68]
  assign _T_2 = io_in_bits_wraddr == 3'h1; // @[ConfigurationMemory.scala 75:65]
  assign _T_4 = io_in_bits_wraddr == 3'h2; // @[ConfigurationMemory.scala 86:63]
  assign _T_6 = io_in_bits_wraddr == 3'h3; // @[ConfigurationMemory.scala 98:66]
  assign _T_8 = io_in_bits_wraddr == 3'h4; // @[ConfigurationMemory.scala 104:29]
  assign _T_9 = io_in_valid & _T_8; // @[ConfigurationMemory.scala 104:20]
  assign _T_10 = $unsigned(io_in_bits_wrdata); // @[ConfigurationMemory.scala 104:90]
  assign _T_11 = _T_10[0]; // @[ConfigurationMemory.scala 104:92]
  assign io_out_bits_confneuralNetsweightMatrix_0_0 = neuralNetsweightMatrixMemory_io_out_bits_0_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_0_1 = neuralNetsweightMatrixMemory_io_out_bits_0_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_0_2 = neuralNetsweightMatrixMemory_io_out_bits_0_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_0_3 = neuralNetsweightMatrixMemory_io_out_bits_0_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_1_0 = neuralNetsweightMatrixMemory_io_out_bits_1_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_1_1 = neuralNetsweightMatrixMemory_io_out_bits_1_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_1_2 = neuralNetsweightMatrixMemory_io_out_bits_1_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_1_3 = neuralNetsweightMatrixMemory_io_out_bits_1_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_2_0 = neuralNetsweightMatrixMemory_io_out_bits_2_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_2_1 = neuralNetsweightMatrixMemory_io_out_bits_2_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_2_2 = neuralNetsweightMatrixMemory_io_out_bits_2_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_2_3 = neuralNetsweightMatrixMemory_io_out_bits_2_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_3_0 = neuralNetsweightMatrixMemory_io_out_bits_3_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_3_1 = neuralNetsweightMatrixMemory_io_out_bits_3_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_3_2 = neuralNetsweightMatrixMemory_io_out_bits_3_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_3_3 = neuralNetsweightMatrixMemory_io_out_bits_3_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_4_0 = neuralNetsweightMatrixMemory_io_out_bits_4_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_4_1 = neuralNetsweightMatrixMemory_io_out_bits_4_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_4_2 = neuralNetsweightMatrixMemory_io_out_bits_4_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_4_3 = neuralNetsweightMatrixMemory_io_out_bits_4_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_5_0 = neuralNetsweightMatrixMemory_io_out_bits_5_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_5_1 = neuralNetsweightMatrixMemory_io_out_bits_5_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_5_2 = neuralNetsweightMatrixMemory_io_out_bits_5_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_5_3 = neuralNetsweightMatrixMemory_io_out_bits_5_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_6_0 = neuralNetsweightMatrixMemory_io_out_bits_6_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_6_1 = neuralNetsweightMatrixMemory_io_out_bits_6_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_6_2 = neuralNetsweightMatrixMemory_io_out_bits_6_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_6_3 = neuralNetsweightMatrixMemory_io_out_bits_6_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_7_0 = neuralNetsweightMatrixMemory_io_out_bits_7_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_7_1 = neuralNetsweightMatrixMemory_io_out_bits_7_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_7_2 = neuralNetsweightMatrixMemory_io_out_bits_7_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_7_3 = neuralNetsweightMatrixMemory_io_out_bits_7_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_8_0 = neuralNetsweightMatrixMemory_io_out_bits_8_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_8_1 = neuralNetsweightMatrixMemory_io_out_bits_8_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_8_2 = neuralNetsweightMatrixMemory_io_out_bits_8_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_8_3 = neuralNetsweightMatrixMemory_io_out_bits_8_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_9_0 = neuralNetsweightMatrixMemory_io_out_bits_9_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_9_1 = neuralNetsweightMatrixMemory_io_out_bits_9_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_9_2 = neuralNetsweightMatrixMemory_io_out_bits_9_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_9_3 = neuralNetsweightMatrixMemory_io_out_bits_9_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_10_0 = neuralNetsweightMatrixMemory_io_out_bits_10_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_10_1 = neuralNetsweightMatrixMemory_io_out_bits_10_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_10_2 = neuralNetsweightMatrixMemory_io_out_bits_10_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_10_3 = neuralNetsweightMatrixMemory_io_out_bits_10_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_11_0 = neuralNetsweightMatrixMemory_io_out_bits_11_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_11_1 = neuralNetsweightMatrixMemory_io_out_bits_11_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_11_2 = neuralNetsweightMatrixMemory_io_out_bits_11_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_11_3 = neuralNetsweightMatrixMemory_io_out_bits_11_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_12_0 = neuralNetsweightMatrixMemory_io_out_bits_12_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_12_1 = neuralNetsweightMatrixMemory_io_out_bits_12_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_12_2 = neuralNetsweightMatrixMemory_io_out_bits_12_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_12_3 = neuralNetsweightMatrixMemory_io_out_bits_12_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_13_0 = neuralNetsweightMatrixMemory_io_out_bits_13_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_13_1 = neuralNetsweightMatrixMemory_io_out_bits_13_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_13_2 = neuralNetsweightMatrixMemory_io_out_bits_13_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_13_3 = neuralNetsweightMatrixMemory_io_out_bits_13_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_14_0 = neuralNetsweightMatrixMemory_io_out_bits_14_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_14_1 = neuralNetsweightMatrixMemory_io_out_bits_14_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_14_2 = neuralNetsweightMatrixMemory_io_out_bits_14_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_14_3 = neuralNetsweightMatrixMemory_io_out_bits_14_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_15_0 = neuralNetsweightMatrixMemory_io_out_bits_15_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_15_1 = neuralNetsweightMatrixMemory_io_out_bits_15_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_15_2 = neuralNetsweightMatrixMemory_io_out_bits_15_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_15_3 = neuralNetsweightMatrixMemory_io_out_bits_15_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_16_0 = neuralNetsweightMatrixMemory_io_out_bits_16_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_16_1 = neuralNetsweightMatrixMemory_io_out_bits_16_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_16_2 = neuralNetsweightMatrixMemory_io_out_bits_16_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_16_3 = neuralNetsweightMatrixMemory_io_out_bits_16_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_17_0 = neuralNetsweightMatrixMemory_io_out_bits_17_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_17_1 = neuralNetsweightMatrixMemory_io_out_bits_17_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_17_2 = neuralNetsweightMatrixMemory_io_out_bits_17_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_17_3 = neuralNetsweightMatrixMemory_io_out_bits_17_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_18_0 = neuralNetsweightMatrixMemory_io_out_bits_18_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_18_1 = neuralNetsweightMatrixMemory_io_out_bits_18_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_18_2 = neuralNetsweightMatrixMemory_io_out_bits_18_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_18_3 = neuralNetsweightMatrixMemory_io_out_bits_18_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_19_0 = neuralNetsweightMatrixMemory_io_out_bits_19_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_19_1 = neuralNetsweightMatrixMemory_io_out_bits_19_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_19_2 = neuralNetsweightMatrixMemory_io_out_bits_19_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_19_3 = neuralNetsweightMatrixMemory_io_out_bits_19_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_20_0 = neuralNetsweightMatrixMemory_io_out_bits_20_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_20_1 = neuralNetsweightMatrixMemory_io_out_bits_20_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_20_2 = neuralNetsweightMatrixMemory_io_out_bits_20_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_20_3 = neuralNetsweightMatrixMemory_io_out_bits_20_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_21_0 = neuralNetsweightMatrixMemory_io_out_bits_21_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_21_1 = neuralNetsweightMatrixMemory_io_out_bits_21_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_21_2 = neuralNetsweightMatrixMemory_io_out_bits_21_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_21_3 = neuralNetsweightMatrixMemory_io_out_bits_21_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_22_0 = neuralNetsweightMatrixMemory_io_out_bits_22_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_22_1 = neuralNetsweightMatrixMemory_io_out_bits_22_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_22_2 = neuralNetsweightMatrixMemory_io_out_bits_22_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_22_3 = neuralNetsweightMatrixMemory_io_out_bits_22_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_23_0 = neuralNetsweightMatrixMemory_io_out_bits_23_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_23_1 = neuralNetsweightMatrixMemory_io_out_bits_23_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_23_2 = neuralNetsweightMatrixMemory_io_out_bits_23_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_23_3 = neuralNetsweightMatrixMemory_io_out_bits_23_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_24_0 = neuralNetsweightMatrixMemory_io_out_bits_24_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_24_1 = neuralNetsweightMatrixMemory_io_out_bits_24_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_24_2 = neuralNetsweightMatrixMemory_io_out_bits_24_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_24_3 = neuralNetsweightMatrixMemory_io_out_bits_24_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_25_0 = neuralNetsweightMatrixMemory_io_out_bits_25_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_25_1 = neuralNetsweightMatrixMemory_io_out_bits_25_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_25_2 = neuralNetsweightMatrixMemory_io_out_bits_25_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_25_3 = neuralNetsweightMatrixMemory_io_out_bits_25_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_26_0 = neuralNetsweightMatrixMemory_io_out_bits_26_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_26_1 = neuralNetsweightMatrixMemory_io_out_bits_26_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_26_2 = neuralNetsweightMatrixMemory_io_out_bits_26_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_26_3 = neuralNetsweightMatrixMemory_io_out_bits_26_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_27_0 = neuralNetsweightMatrixMemory_io_out_bits_27_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_27_1 = neuralNetsweightMatrixMemory_io_out_bits_27_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_27_2 = neuralNetsweightMatrixMemory_io_out_bits_27_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_27_3 = neuralNetsweightMatrixMemory_io_out_bits_27_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_28_0 = neuralNetsweightMatrixMemory_io_out_bits_28_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_28_1 = neuralNetsweightMatrixMemory_io_out_bits_28_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_28_2 = neuralNetsweightMatrixMemory_io_out_bits_28_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_28_3 = neuralNetsweightMatrixMemory_io_out_bits_28_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_29_0 = neuralNetsweightMatrixMemory_io_out_bits_29_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_29_1 = neuralNetsweightMatrixMemory_io_out_bits_29_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_29_2 = neuralNetsweightMatrixMemory_io_out_bits_29_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_29_3 = neuralNetsweightMatrixMemory_io_out_bits_29_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_30_0 = neuralNetsweightMatrixMemory_io_out_bits_30_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_30_1 = neuralNetsweightMatrixMemory_io_out_bits_30_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_30_2 = neuralNetsweightMatrixMemory_io_out_bits_30_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_30_3 = neuralNetsweightMatrixMemory_io_out_bits_30_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_31_0 = neuralNetsweightMatrixMemory_io_out_bits_31_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_31_1 = neuralNetsweightMatrixMemory_io_out_bits_31_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_31_2 = neuralNetsweightMatrixMemory_io_out_bits_31_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_31_3 = neuralNetsweightMatrixMemory_io_out_bits_31_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_32_0 = neuralNetsweightMatrixMemory_io_out_bits_32_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_32_1 = neuralNetsweightMatrixMemory_io_out_bits_32_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_32_2 = neuralNetsweightMatrixMemory_io_out_bits_32_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_32_3 = neuralNetsweightMatrixMemory_io_out_bits_32_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_33_0 = neuralNetsweightMatrixMemory_io_out_bits_33_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_33_1 = neuralNetsweightMatrixMemory_io_out_bits_33_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_33_2 = neuralNetsweightMatrixMemory_io_out_bits_33_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_33_3 = neuralNetsweightMatrixMemory_io_out_bits_33_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_34_0 = neuralNetsweightMatrixMemory_io_out_bits_34_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_34_1 = neuralNetsweightMatrixMemory_io_out_bits_34_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_34_2 = neuralNetsweightMatrixMemory_io_out_bits_34_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_34_3 = neuralNetsweightMatrixMemory_io_out_bits_34_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_35_0 = neuralNetsweightMatrixMemory_io_out_bits_35_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_35_1 = neuralNetsweightMatrixMemory_io_out_bits_35_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_35_2 = neuralNetsweightMatrixMemory_io_out_bits_35_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_35_3 = neuralNetsweightMatrixMemory_io_out_bits_35_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_36_0 = neuralNetsweightMatrixMemory_io_out_bits_36_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_36_1 = neuralNetsweightMatrixMemory_io_out_bits_36_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_36_2 = neuralNetsweightMatrixMemory_io_out_bits_36_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_36_3 = neuralNetsweightMatrixMemory_io_out_bits_36_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_37_0 = neuralNetsweightMatrixMemory_io_out_bits_37_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_37_1 = neuralNetsweightMatrixMemory_io_out_bits_37_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_37_2 = neuralNetsweightMatrixMemory_io_out_bits_37_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_37_3 = neuralNetsweightMatrixMemory_io_out_bits_37_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_38_0 = neuralNetsweightMatrixMemory_io_out_bits_38_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_38_1 = neuralNetsweightMatrixMemory_io_out_bits_38_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_38_2 = neuralNetsweightMatrixMemory_io_out_bits_38_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_38_3 = neuralNetsweightMatrixMemory_io_out_bits_38_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_39_0 = neuralNetsweightMatrixMemory_io_out_bits_39_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_39_1 = neuralNetsweightMatrixMemory_io_out_bits_39_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_39_2 = neuralNetsweightMatrixMemory_io_out_bits_39_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_39_3 = neuralNetsweightMatrixMemory_io_out_bits_39_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_40_0 = neuralNetsweightMatrixMemory_io_out_bits_40_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_40_1 = neuralNetsweightMatrixMemory_io_out_bits_40_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_40_2 = neuralNetsweightMatrixMemory_io_out_bits_40_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_40_3 = neuralNetsweightMatrixMemory_io_out_bits_40_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_41_0 = neuralNetsweightMatrixMemory_io_out_bits_41_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_41_1 = neuralNetsweightMatrixMemory_io_out_bits_41_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_41_2 = neuralNetsweightMatrixMemory_io_out_bits_41_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_41_3 = neuralNetsweightMatrixMemory_io_out_bits_41_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_42_0 = neuralNetsweightMatrixMemory_io_out_bits_42_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_42_1 = neuralNetsweightMatrixMemory_io_out_bits_42_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_42_2 = neuralNetsweightMatrixMemory_io_out_bits_42_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_42_3 = neuralNetsweightMatrixMemory_io_out_bits_42_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_43_0 = neuralNetsweightMatrixMemory_io_out_bits_43_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_43_1 = neuralNetsweightMatrixMemory_io_out_bits_43_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_43_2 = neuralNetsweightMatrixMemory_io_out_bits_43_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_43_3 = neuralNetsweightMatrixMemory_io_out_bits_43_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_44_0 = neuralNetsweightMatrixMemory_io_out_bits_44_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_44_1 = neuralNetsweightMatrixMemory_io_out_bits_44_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_44_2 = neuralNetsweightMatrixMemory_io_out_bits_44_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_44_3 = neuralNetsweightMatrixMemory_io_out_bits_44_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_45_0 = neuralNetsweightMatrixMemory_io_out_bits_45_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_45_1 = neuralNetsweightMatrixMemory_io_out_bits_45_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_45_2 = neuralNetsweightMatrixMemory_io_out_bits_45_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_45_3 = neuralNetsweightMatrixMemory_io_out_bits_45_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_46_0 = neuralNetsweightMatrixMemory_io_out_bits_46_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_46_1 = neuralNetsweightMatrixMemory_io_out_bits_46_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_46_2 = neuralNetsweightMatrixMemory_io_out_bits_46_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_46_3 = neuralNetsweightMatrixMemory_io_out_bits_46_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_47_0 = neuralNetsweightMatrixMemory_io_out_bits_47_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_47_1 = neuralNetsweightMatrixMemory_io_out_bits_47_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_47_2 = neuralNetsweightMatrixMemory_io_out_bits_47_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_47_3 = neuralNetsweightMatrixMemory_io_out_bits_47_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_48_0 = neuralNetsweightMatrixMemory_io_out_bits_48_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_48_1 = neuralNetsweightMatrixMemory_io_out_bits_48_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_48_2 = neuralNetsweightMatrixMemory_io_out_bits_48_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_48_3 = neuralNetsweightMatrixMemory_io_out_bits_48_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_49_0 = neuralNetsweightMatrixMemory_io_out_bits_49_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_49_1 = neuralNetsweightMatrixMemory_io_out_bits_49_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_49_2 = neuralNetsweightMatrixMemory_io_out_bits_49_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_49_3 = neuralNetsweightMatrixMemory_io_out_bits_49_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_50_0 = neuralNetsweightMatrixMemory_io_out_bits_50_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_50_1 = neuralNetsweightMatrixMemory_io_out_bits_50_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_50_2 = neuralNetsweightMatrixMemory_io_out_bits_50_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_50_3 = neuralNetsweightMatrixMemory_io_out_bits_50_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_51_0 = neuralNetsweightMatrixMemory_io_out_bits_51_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_51_1 = neuralNetsweightMatrixMemory_io_out_bits_51_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_51_2 = neuralNetsweightMatrixMemory_io_out_bits_51_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_51_3 = neuralNetsweightMatrixMemory_io_out_bits_51_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_52_0 = neuralNetsweightMatrixMemory_io_out_bits_52_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_52_1 = neuralNetsweightMatrixMemory_io_out_bits_52_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_52_2 = neuralNetsweightMatrixMemory_io_out_bits_52_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_52_3 = neuralNetsweightMatrixMemory_io_out_bits_52_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_53_0 = neuralNetsweightMatrixMemory_io_out_bits_53_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_53_1 = neuralNetsweightMatrixMemory_io_out_bits_53_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_53_2 = neuralNetsweightMatrixMemory_io_out_bits_53_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_53_3 = neuralNetsweightMatrixMemory_io_out_bits_53_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_54_0 = neuralNetsweightMatrixMemory_io_out_bits_54_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_54_1 = neuralNetsweightMatrixMemory_io_out_bits_54_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_54_2 = neuralNetsweightMatrixMemory_io_out_bits_54_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_54_3 = neuralNetsweightMatrixMemory_io_out_bits_54_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_55_0 = neuralNetsweightMatrixMemory_io_out_bits_55_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_55_1 = neuralNetsweightMatrixMemory_io_out_bits_55_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_55_2 = neuralNetsweightMatrixMemory_io_out_bits_55_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_55_3 = neuralNetsweightMatrixMemory_io_out_bits_55_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_56_0 = neuralNetsweightMatrixMemory_io_out_bits_56_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_56_1 = neuralNetsweightMatrixMemory_io_out_bits_56_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_56_2 = neuralNetsweightMatrixMemory_io_out_bits_56_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_56_3 = neuralNetsweightMatrixMemory_io_out_bits_56_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_57_0 = neuralNetsweightMatrixMemory_io_out_bits_57_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_57_1 = neuralNetsweightMatrixMemory_io_out_bits_57_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_57_2 = neuralNetsweightMatrixMemory_io_out_bits_57_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_57_3 = neuralNetsweightMatrixMemory_io_out_bits_57_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_58_0 = neuralNetsweightMatrixMemory_io_out_bits_58_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_58_1 = neuralNetsweightMatrixMemory_io_out_bits_58_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_58_2 = neuralNetsweightMatrixMemory_io_out_bits_58_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_58_3 = neuralNetsweightMatrixMemory_io_out_bits_58_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_59_0 = neuralNetsweightMatrixMemory_io_out_bits_59_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_59_1 = neuralNetsweightMatrixMemory_io_out_bits_59_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_59_2 = neuralNetsweightMatrixMemory_io_out_bits_59_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_59_3 = neuralNetsweightMatrixMemory_io_out_bits_59_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_60_0 = neuralNetsweightMatrixMemory_io_out_bits_60_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_60_1 = neuralNetsweightMatrixMemory_io_out_bits_60_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_60_2 = neuralNetsweightMatrixMemory_io_out_bits_60_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_60_3 = neuralNetsweightMatrixMemory_io_out_bits_60_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_61_0 = neuralNetsweightMatrixMemory_io_out_bits_61_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_61_1 = neuralNetsweightMatrixMemory_io_out_bits_61_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_61_2 = neuralNetsweightMatrixMemory_io_out_bits_61_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_61_3 = neuralNetsweightMatrixMemory_io_out_bits_61_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_62_0 = neuralNetsweightMatrixMemory_io_out_bits_62_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_62_1 = neuralNetsweightMatrixMemory_io_out_bits_62_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_62_2 = neuralNetsweightMatrixMemory_io_out_bits_62_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_62_3 = neuralNetsweightMatrixMemory_io_out_bits_62_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_63_0 = neuralNetsweightMatrixMemory_io_out_bits_63_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_63_1 = neuralNetsweightMatrixMemory_io_out_bits_63_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_63_2 = neuralNetsweightMatrixMemory_io_out_bits_63_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_63_3 = neuralNetsweightMatrixMemory_io_out_bits_63_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_64_0 = neuralNetsweightMatrixMemory_io_out_bits_64_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_64_1 = neuralNetsweightMatrixMemory_io_out_bits_64_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_64_2 = neuralNetsweightMatrixMemory_io_out_bits_64_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_64_3 = neuralNetsweightMatrixMemory_io_out_bits_64_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_65_0 = neuralNetsweightMatrixMemory_io_out_bits_65_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_65_1 = neuralNetsweightMatrixMemory_io_out_bits_65_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_65_2 = neuralNetsweightMatrixMemory_io_out_bits_65_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_65_3 = neuralNetsweightMatrixMemory_io_out_bits_65_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_66_0 = neuralNetsweightMatrixMemory_io_out_bits_66_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_66_1 = neuralNetsweightMatrixMemory_io_out_bits_66_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_66_2 = neuralNetsweightMatrixMemory_io_out_bits_66_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_66_3 = neuralNetsweightMatrixMemory_io_out_bits_66_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_67_0 = neuralNetsweightMatrixMemory_io_out_bits_67_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_67_1 = neuralNetsweightMatrixMemory_io_out_bits_67_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_67_2 = neuralNetsweightMatrixMemory_io_out_bits_67_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_67_3 = neuralNetsweightMatrixMemory_io_out_bits_67_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_68_0 = neuralNetsweightMatrixMemory_io_out_bits_68_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_68_1 = neuralNetsweightMatrixMemory_io_out_bits_68_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_68_2 = neuralNetsweightMatrixMemory_io_out_bits_68_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_68_3 = neuralNetsweightMatrixMemory_io_out_bits_68_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_69_0 = neuralNetsweightMatrixMemory_io_out_bits_69_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_69_1 = neuralNetsweightMatrixMemory_io_out_bits_69_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_69_2 = neuralNetsweightMatrixMemory_io_out_bits_69_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_69_3 = neuralNetsweightMatrixMemory_io_out_bits_69_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_70_0 = neuralNetsweightMatrixMemory_io_out_bits_70_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_70_1 = neuralNetsweightMatrixMemory_io_out_bits_70_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_70_2 = neuralNetsweightMatrixMemory_io_out_bits_70_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_70_3 = neuralNetsweightMatrixMemory_io_out_bits_70_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_71_0 = neuralNetsweightMatrixMemory_io_out_bits_71_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_71_1 = neuralNetsweightMatrixMemory_io_out_bits_71_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_71_2 = neuralNetsweightMatrixMemory_io_out_bits_71_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_71_3 = neuralNetsweightMatrixMemory_io_out_bits_71_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_72_0 = neuralNetsweightMatrixMemory_io_out_bits_72_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_72_1 = neuralNetsweightMatrixMemory_io_out_bits_72_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_72_2 = neuralNetsweightMatrixMemory_io_out_bits_72_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_72_3 = neuralNetsweightMatrixMemory_io_out_bits_72_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_73_0 = neuralNetsweightMatrixMemory_io_out_bits_73_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_73_1 = neuralNetsweightMatrixMemory_io_out_bits_73_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_73_2 = neuralNetsweightMatrixMemory_io_out_bits_73_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_73_3 = neuralNetsweightMatrixMemory_io_out_bits_73_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_74_0 = neuralNetsweightMatrixMemory_io_out_bits_74_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_74_1 = neuralNetsweightMatrixMemory_io_out_bits_74_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_74_2 = neuralNetsweightMatrixMemory_io_out_bits_74_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_74_3 = neuralNetsweightMatrixMemory_io_out_bits_74_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_75_0 = neuralNetsweightMatrixMemory_io_out_bits_75_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_75_1 = neuralNetsweightMatrixMemory_io_out_bits_75_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_75_2 = neuralNetsweightMatrixMemory_io_out_bits_75_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_75_3 = neuralNetsweightMatrixMemory_io_out_bits_75_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_76_0 = neuralNetsweightMatrixMemory_io_out_bits_76_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_76_1 = neuralNetsweightMatrixMemory_io_out_bits_76_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_76_2 = neuralNetsweightMatrixMemory_io_out_bits_76_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_76_3 = neuralNetsweightMatrixMemory_io_out_bits_76_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_77_0 = neuralNetsweightMatrixMemory_io_out_bits_77_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_77_1 = neuralNetsweightMatrixMemory_io_out_bits_77_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_77_2 = neuralNetsweightMatrixMemory_io_out_bits_77_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_77_3 = neuralNetsweightMatrixMemory_io_out_bits_77_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_78_0 = neuralNetsweightMatrixMemory_io_out_bits_78_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_78_1 = neuralNetsweightMatrixMemory_io_out_bits_78_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_78_2 = neuralNetsweightMatrixMemory_io_out_bits_78_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_78_3 = neuralNetsweightMatrixMemory_io_out_bits_78_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_79_0 = neuralNetsweightMatrixMemory_io_out_bits_79_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_79_1 = neuralNetsweightMatrixMemory_io_out_bits_79_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_79_2 = neuralNetsweightMatrixMemory_io_out_bits_79_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_79_3 = neuralNetsweightMatrixMemory_io_out_bits_79_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_80_0 = neuralNetsweightMatrixMemory_io_out_bits_80_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_80_1 = neuralNetsweightMatrixMemory_io_out_bits_80_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_80_2 = neuralNetsweightMatrixMemory_io_out_bits_80_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_80_3 = neuralNetsweightMatrixMemory_io_out_bits_80_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_81_0 = neuralNetsweightMatrixMemory_io_out_bits_81_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_81_1 = neuralNetsweightMatrixMemory_io_out_bits_81_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_81_2 = neuralNetsweightMatrixMemory_io_out_bits_81_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_81_3 = neuralNetsweightMatrixMemory_io_out_bits_81_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_82_0 = neuralNetsweightMatrixMemory_io_out_bits_82_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_82_1 = neuralNetsweightMatrixMemory_io_out_bits_82_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_82_2 = neuralNetsweightMatrixMemory_io_out_bits_82_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_82_3 = neuralNetsweightMatrixMemory_io_out_bits_82_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_83_0 = neuralNetsweightMatrixMemory_io_out_bits_83_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_83_1 = neuralNetsweightMatrixMemory_io_out_bits_83_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_83_2 = neuralNetsweightMatrixMemory_io_out_bits_83_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_83_3 = neuralNetsweightMatrixMemory_io_out_bits_83_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_84_0 = neuralNetsweightMatrixMemory_io_out_bits_84_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_84_1 = neuralNetsweightMatrixMemory_io_out_bits_84_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_84_2 = neuralNetsweightMatrixMemory_io_out_bits_84_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_84_3 = neuralNetsweightMatrixMemory_io_out_bits_84_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_85_0 = neuralNetsweightMatrixMemory_io_out_bits_85_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_85_1 = neuralNetsweightMatrixMemory_io_out_bits_85_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_85_2 = neuralNetsweightMatrixMemory_io_out_bits_85_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_85_3 = neuralNetsweightMatrixMemory_io_out_bits_85_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_86_0 = neuralNetsweightMatrixMemory_io_out_bits_86_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_86_1 = neuralNetsweightMatrixMemory_io_out_bits_86_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_86_2 = neuralNetsweightMatrixMemory_io_out_bits_86_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_86_3 = neuralNetsweightMatrixMemory_io_out_bits_86_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_87_0 = neuralNetsweightMatrixMemory_io_out_bits_87_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_87_1 = neuralNetsweightMatrixMemory_io_out_bits_87_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_87_2 = neuralNetsweightMatrixMemory_io_out_bits_87_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_87_3 = neuralNetsweightMatrixMemory_io_out_bits_87_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_88_0 = neuralNetsweightMatrixMemory_io_out_bits_88_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_88_1 = neuralNetsweightMatrixMemory_io_out_bits_88_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_88_2 = neuralNetsweightMatrixMemory_io_out_bits_88_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_88_3 = neuralNetsweightMatrixMemory_io_out_bits_88_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_89_0 = neuralNetsweightMatrixMemory_io_out_bits_89_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_89_1 = neuralNetsweightMatrixMemory_io_out_bits_89_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_89_2 = neuralNetsweightMatrixMemory_io_out_bits_89_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_89_3 = neuralNetsweightMatrixMemory_io_out_bits_89_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_90_0 = neuralNetsweightMatrixMemory_io_out_bits_90_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_90_1 = neuralNetsweightMatrixMemory_io_out_bits_90_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_90_2 = neuralNetsweightMatrixMemory_io_out_bits_90_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_90_3 = neuralNetsweightMatrixMemory_io_out_bits_90_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_91_0 = neuralNetsweightMatrixMemory_io_out_bits_91_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_91_1 = neuralNetsweightMatrixMemory_io_out_bits_91_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_91_2 = neuralNetsweightMatrixMemory_io_out_bits_91_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_91_3 = neuralNetsweightMatrixMemory_io_out_bits_91_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_92_0 = neuralNetsweightMatrixMemory_io_out_bits_92_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_92_1 = neuralNetsweightMatrixMemory_io_out_bits_92_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_92_2 = neuralNetsweightMatrixMemory_io_out_bits_92_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_92_3 = neuralNetsweightMatrixMemory_io_out_bits_92_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_93_0 = neuralNetsweightMatrixMemory_io_out_bits_93_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_93_1 = neuralNetsweightMatrixMemory_io_out_bits_93_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_93_2 = neuralNetsweightMatrixMemory_io_out_bits_93_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_93_3 = neuralNetsweightMatrixMemory_io_out_bits_93_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_94_0 = neuralNetsweightMatrixMemory_io_out_bits_94_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_94_1 = neuralNetsweightMatrixMemory_io_out_bits_94_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_94_2 = neuralNetsweightMatrixMemory_io_out_bits_94_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_94_3 = neuralNetsweightMatrixMemory_io_out_bits_94_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_95_0 = neuralNetsweightMatrixMemory_io_out_bits_95_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_95_1 = neuralNetsweightMatrixMemory_io_out_bits_95_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_95_2 = neuralNetsweightMatrixMemory_io_out_bits_95_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_95_3 = neuralNetsweightMatrixMemory_io_out_bits_95_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_96_0 = neuralNetsweightMatrixMemory_io_out_bits_96_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_96_1 = neuralNetsweightMatrixMemory_io_out_bits_96_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_96_2 = neuralNetsweightMatrixMemory_io_out_bits_96_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_96_3 = neuralNetsweightMatrixMemory_io_out_bits_96_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_97_0 = neuralNetsweightMatrixMemory_io_out_bits_97_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_97_1 = neuralNetsweightMatrixMemory_io_out_bits_97_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_97_2 = neuralNetsweightMatrixMemory_io_out_bits_97_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_97_3 = neuralNetsweightMatrixMemory_io_out_bits_97_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_98_0 = neuralNetsweightMatrixMemory_io_out_bits_98_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_98_1 = neuralNetsweightMatrixMemory_io_out_bits_98_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_98_2 = neuralNetsweightMatrixMemory_io_out_bits_98_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_98_3 = neuralNetsweightMatrixMemory_io_out_bits_98_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_99_0 = neuralNetsweightMatrixMemory_io_out_bits_99_0; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_99_1 = neuralNetsweightMatrixMemory_io_out_bits_99_1; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_99_2 = neuralNetsweightMatrixMemory_io_out_bits_99_2; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightMatrix_99_3 = neuralNetsweightMatrixMemory_io_out_bits_99_3; // @[ConfigurationMemory.scala 64:42]
  assign io_out_bits_confneuralNetsweightVec_0 = neuralNetsweightVecMemory_io_out_bits_0_0; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_1 = neuralNetsweightVecMemory_io_out_bits_0_1; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_2 = neuralNetsweightVecMemory_io_out_bits_0_2; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_3 = neuralNetsweightVecMemory_io_out_bits_0_3; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_4 = neuralNetsweightVecMemory_io_out_bits_0_4; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_5 = neuralNetsweightVecMemory_io_out_bits_0_5; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_6 = neuralNetsweightVecMemory_io_out_bits_0_6; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_7 = neuralNetsweightVecMemory_io_out_bits_0_7; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_8 = neuralNetsweightVecMemory_io_out_bits_0_8; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_9 = neuralNetsweightVecMemory_io_out_bits_0_9; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_10 = neuralNetsweightVecMemory_io_out_bits_0_10; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_11 = neuralNetsweightVecMemory_io_out_bits_0_11; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_12 = neuralNetsweightVecMemory_io_out_bits_0_12; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_13 = neuralNetsweightVecMemory_io_out_bits_0_13; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_14 = neuralNetsweightVecMemory_io_out_bits_0_14; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_15 = neuralNetsweightVecMemory_io_out_bits_0_15; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_16 = neuralNetsweightVecMemory_io_out_bits_0_16; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_17 = neuralNetsweightVecMemory_io_out_bits_0_17; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_18 = neuralNetsweightVecMemory_io_out_bits_0_18; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_19 = neuralNetsweightVecMemory_io_out_bits_0_19; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_20 = neuralNetsweightVecMemory_io_out_bits_0_20; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_21 = neuralNetsweightVecMemory_io_out_bits_0_21; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_22 = neuralNetsweightVecMemory_io_out_bits_0_22; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_23 = neuralNetsweightVecMemory_io_out_bits_0_23; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_24 = neuralNetsweightVecMemory_io_out_bits_0_24; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_25 = neuralNetsweightVecMemory_io_out_bits_0_25; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_26 = neuralNetsweightVecMemory_io_out_bits_0_26; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_27 = neuralNetsweightVecMemory_io_out_bits_0_27; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_28 = neuralNetsweightVecMemory_io_out_bits_0_28; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_29 = neuralNetsweightVecMemory_io_out_bits_0_29; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_30 = neuralNetsweightVecMemory_io_out_bits_0_30; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_31 = neuralNetsweightVecMemory_io_out_bits_0_31; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_32 = neuralNetsweightVecMemory_io_out_bits_0_32; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_33 = neuralNetsweightVecMemory_io_out_bits_0_33; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_34 = neuralNetsweightVecMemory_io_out_bits_0_34; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_35 = neuralNetsweightVecMemory_io_out_bits_0_35; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_36 = neuralNetsweightVecMemory_io_out_bits_0_36; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_37 = neuralNetsweightVecMemory_io_out_bits_0_37; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_38 = neuralNetsweightVecMemory_io_out_bits_0_38; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_39 = neuralNetsweightVecMemory_io_out_bits_0_39; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_40 = neuralNetsweightVecMemory_io_out_bits_0_40; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_41 = neuralNetsweightVecMemory_io_out_bits_0_41; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_42 = neuralNetsweightVecMemory_io_out_bits_0_42; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_43 = neuralNetsweightVecMemory_io_out_bits_0_43; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_44 = neuralNetsweightVecMemory_io_out_bits_0_44; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_45 = neuralNetsweightVecMemory_io_out_bits_0_45; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_46 = neuralNetsweightVecMemory_io_out_bits_0_46; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_47 = neuralNetsweightVecMemory_io_out_bits_0_47; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_48 = neuralNetsweightVecMemory_io_out_bits_0_48; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_49 = neuralNetsweightVecMemory_io_out_bits_0_49; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_50 = neuralNetsweightVecMemory_io_out_bits_0_50; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_51 = neuralNetsweightVecMemory_io_out_bits_0_51; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_52 = neuralNetsweightVecMemory_io_out_bits_0_52; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_53 = neuralNetsweightVecMemory_io_out_bits_0_53; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_54 = neuralNetsweightVecMemory_io_out_bits_0_54; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_55 = neuralNetsweightVecMemory_io_out_bits_0_55; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_56 = neuralNetsweightVecMemory_io_out_bits_0_56; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_57 = neuralNetsweightVecMemory_io_out_bits_0_57; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_58 = neuralNetsweightVecMemory_io_out_bits_0_58; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_59 = neuralNetsweightVecMemory_io_out_bits_0_59; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_60 = neuralNetsweightVecMemory_io_out_bits_0_60; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_61 = neuralNetsweightVecMemory_io_out_bits_0_61; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_62 = neuralNetsweightVecMemory_io_out_bits_0_62; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_63 = neuralNetsweightVecMemory_io_out_bits_0_63; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_64 = neuralNetsweightVecMemory_io_out_bits_0_64; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_65 = neuralNetsweightVecMemory_io_out_bits_0_65; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_66 = neuralNetsweightVecMemory_io_out_bits_0_66; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_67 = neuralNetsweightVecMemory_io_out_bits_0_67; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_68 = neuralNetsweightVecMemory_io_out_bits_0_68; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_69 = neuralNetsweightVecMemory_io_out_bits_0_69; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_70 = neuralNetsweightVecMemory_io_out_bits_0_70; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_71 = neuralNetsweightVecMemory_io_out_bits_0_71; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_72 = neuralNetsweightVecMemory_io_out_bits_0_72; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_73 = neuralNetsweightVecMemory_io_out_bits_0_73; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_74 = neuralNetsweightVecMemory_io_out_bits_0_74; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_75 = neuralNetsweightVecMemory_io_out_bits_0_75; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_76 = neuralNetsweightVecMemory_io_out_bits_0_76; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_77 = neuralNetsweightVecMemory_io_out_bits_0_77; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_78 = neuralNetsweightVecMemory_io_out_bits_0_78; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_79 = neuralNetsweightVecMemory_io_out_bits_0_79; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_80 = neuralNetsweightVecMemory_io_out_bits_0_80; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_81 = neuralNetsweightVecMemory_io_out_bits_0_81; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_82 = neuralNetsweightVecMemory_io_out_bits_0_82; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_83 = neuralNetsweightVecMemory_io_out_bits_0_83; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_84 = neuralNetsweightVecMemory_io_out_bits_0_84; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_85 = neuralNetsweightVecMemory_io_out_bits_0_85; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_86 = neuralNetsweightVecMemory_io_out_bits_0_86; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_87 = neuralNetsweightVecMemory_io_out_bits_0_87; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_88 = neuralNetsweightVecMemory_io_out_bits_0_88; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_89 = neuralNetsweightVecMemory_io_out_bits_0_89; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_90 = neuralNetsweightVecMemory_io_out_bits_0_90; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_91 = neuralNetsweightVecMemory_io_out_bits_0_91; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_92 = neuralNetsweightVecMemory_io_out_bits_0_92; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_93 = neuralNetsweightVecMemory_io_out_bits_0_93; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_94 = neuralNetsweightVecMemory_io_out_bits_0_94; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_95 = neuralNetsweightVecMemory_io_out_bits_0_95; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_96 = neuralNetsweightVecMemory_io_out_bits_0_96; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_97 = neuralNetsweightVecMemory_io_out_bits_0_97; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_98 = neuralNetsweightVecMemory_io_out_bits_0_98; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsweightVec_99 = neuralNetsweightVecMemory_io_out_bits_0_99; // @[ConfigurationMemory.scala 76:39]
  assign io_out_bits_confneuralNetsbiasVec_0 = neuralNetsbiasVecMemory_io_out_bits_0_0; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_1 = neuralNetsbiasVecMemory_io_out_bits_0_1; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_2 = neuralNetsbiasVecMemory_io_out_bits_0_2; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_3 = neuralNetsbiasVecMemory_io_out_bits_0_3; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_4 = neuralNetsbiasVecMemory_io_out_bits_0_4; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_5 = neuralNetsbiasVecMemory_io_out_bits_0_5; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_6 = neuralNetsbiasVecMemory_io_out_bits_0_6; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_7 = neuralNetsbiasVecMemory_io_out_bits_0_7; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_8 = neuralNetsbiasVecMemory_io_out_bits_0_8; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_9 = neuralNetsbiasVecMemory_io_out_bits_0_9; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_10 = neuralNetsbiasVecMemory_io_out_bits_0_10; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_11 = neuralNetsbiasVecMemory_io_out_bits_0_11; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_12 = neuralNetsbiasVecMemory_io_out_bits_0_12; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_13 = neuralNetsbiasVecMemory_io_out_bits_0_13; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_14 = neuralNetsbiasVecMemory_io_out_bits_0_14; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_15 = neuralNetsbiasVecMemory_io_out_bits_0_15; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_16 = neuralNetsbiasVecMemory_io_out_bits_0_16; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_17 = neuralNetsbiasVecMemory_io_out_bits_0_17; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_18 = neuralNetsbiasVecMemory_io_out_bits_0_18; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_19 = neuralNetsbiasVecMemory_io_out_bits_0_19; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_20 = neuralNetsbiasVecMemory_io_out_bits_0_20; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_21 = neuralNetsbiasVecMemory_io_out_bits_0_21; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_22 = neuralNetsbiasVecMemory_io_out_bits_0_22; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_23 = neuralNetsbiasVecMemory_io_out_bits_0_23; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_24 = neuralNetsbiasVecMemory_io_out_bits_0_24; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_25 = neuralNetsbiasVecMemory_io_out_bits_0_25; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_26 = neuralNetsbiasVecMemory_io_out_bits_0_26; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_27 = neuralNetsbiasVecMemory_io_out_bits_0_27; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_28 = neuralNetsbiasVecMemory_io_out_bits_0_28; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_29 = neuralNetsbiasVecMemory_io_out_bits_0_29; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_30 = neuralNetsbiasVecMemory_io_out_bits_0_30; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_31 = neuralNetsbiasVecMemory_io_out_bits_0_31; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_32 = neuralNetsbiasVecMemory_io_out_bits_0_32; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_33 = neuralNetsbiasVecMemory_io_out_bits_0_33; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_34 = neuralNetsbiasVecMemory_io_out_bits_0_34; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_35 = neuralNetsbiasVecMemory_io_out_bits_0_35; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_36 = neuralNetsbiasVecMemory_io_out_bits_0_36; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_37 = neuralNetsbiasVecMemory_io_out_bits_0_37; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_38 = neuralNetsbiasVecMemory_io_out_bits_0_38; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_39 = neuralNetsbiasVecMemory_io_out_bits_0_39; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_40 = neuralNetsbiasVecMemory_io_out_bits_0_40; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_41 = neuralNetsbiasVecMemory_io_out_bits_0_41; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_42 = neuralNetsbiasVecMemory_io_out_bits_0_42; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_43 = neuralNetsbiasVecMemory_io_out_bits_0_43; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_44 = neuralNetsbiasVecMemory_io_out_bits_0_44; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_45 = neuralNetsbiasVecMemory_io_out_bits_0_45; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_46 = neuralNetsbiasVecMemory_io_out_bits_0_46; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_47 = neuralNetsbiasVecMemory_io_out_bits_0_47; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_48 = neuralNetsbiasVecMemory_io_out_bits_0_48; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_49 = neuralNetsbiasVecMemory_io_out_bits_0_49; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_50 = neuralNetsbiasVecMemory_io_out_bits_0_50; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_51 = neuralNetsbiasVecMemory_io_out_bits_0_51; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_52 = neuralNetsbiasVecMemory_io_out_bits_0_52; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_53 = neuralNetsbiasVecMemory_io_out_bits_0_53; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_54 = neuralNetsbiasVecMemory_io_out_bits_0_54; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_55 = neuralNetsbiasVecMemory_io_out_bits_0_55; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_56 = neuralNetsbiasVecMemory_io_out_bits_0_56; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_57 = neuralNetsbiasVecMemory_io_out_bits_0_57; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_58 = neuralNetsbiasVecMemory_io_out_bits_0_58; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_59 = neuralNetsbiasVecMemory_io_out_bits_0_59; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_60 = neuralNetsbiasVecMemory_io_out_bits_0_60; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_61 = neuralNetsbiasVecMemory_io_out_bits_0_61; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_62 = neuralNetsbiasVecMemory_io_out_bits_0_62; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_63 = neuralNetsbiasVecMemory_io_out_bits_0_63; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_64 = neuralNetsbiasVecMemory_io_out_bits_0_64; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_65 = neuralNetsbiasVecMemory_io_out_bits_0_65; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_66 = neuralNetsbiasVecMemory_io_out_bits_0_66; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_67 = neuralNetsbiasVecMemory_io_out_bits_0_67; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_68 = neuralNetsbiasVecMemory_io_out_bits_0_68; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_69 = neuralNetsbiasVecMemory_io_out_bits_0_69; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_70 = neuralNetsbiasVecMemory_io_out_bits_0_70; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_71 = neuralNetsbiasVecMemory_io_out_bits_0_71; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_72 = neuralNetsbiasVecMemory_io_out_bits_0_72; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_73 = neuralNetsbiasVecMemory_io_out_bits_0_73; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_74 = neuralNetsbiasVecMemory_io_out_bits_0_74; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_75 = neuralNetsbiasVecMemory_io_out_bits_0_75; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_76 = neuralNetsbiasVecMemory_io_out_bits_0_76; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_77 = neuralNetsbiasVecMemory_io_out_bits_0_77; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_78 = neuralNetsbiasVecMemory_io_out_bits_0_78; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_79 = neuralNetsbiasVecMemory_io_out_bits_0_79; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_80 = neuralNetsbiasVecMemory_io_out_bits_0_80; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_81 = neuralNetsbiasVecMemory_io_out_bits_0_81; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_82 = neuralNetsbiasVecMemory_io_out_bits_0_82; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_83 = neuralNetsbiasVecMemory_io_out_bits_0_83; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_84 = neuralNetsbiasVecMemory_io_out_bits_0_84; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_85 = neuralNetsbiasVecMemory_io_out_bits_0_85; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_86 = neuralNetsbiasVecMemory_io_out_bits_0_86; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_87 = neuralNetsbiasVecMemory_io_out_bits_0_87; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_88 = neuralNetsbiasVecMemory_io_out_bits_0_88; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_89 = neuralNetsbiasVecMemory_io_out_bits_0_89; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_90 = neuralNetsbiasVecMemory_io_out_bits_0_90; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_91 = neuralNetsbiasVecMemory_io_out_bits_0_91; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_92 = neuralNetsbiasVecMemory_io_out_bits_0_92; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_93 = neuralNetsbiasVecMemory_io_out_bits_0_93; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_94 = neuralNetsbiasVecMemory_io_out_bits_0_94; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_95 = neuralNetsbiasVecMemory_io_out_bits_0_95; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_96 = neuralNetsbiasVecMemory_io_out_bits_0_96; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_97 = neuralNetsbiasVecMemory_io_out_bits_0_97; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_98 = neuralNetsbiasVecMemory_io_out_bits_0_98; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasVec_99 = neuralNetsbiasVecMemory_io_out_bits_0_99; // @[ConfigurationMemory.scala 87:37]
  assign io_out_bits_confneuralNetsbiasScalar_0 = neuralNetsbiasScalarMemory_io_out_bits_0_0; // @[ConfigurationMemory.scala 99:40]
  assign io_out_bits_confInputMuxSel = inputMuxSel; // @[ConfigurationMemory.scala 105:31]
  assign neuralNetsweightMatrixMemory_clock = clock;
  assign neuralNetsweightMatrixMemory_reset = reset;
  assign neuralNetsweightMatrixMemory_io_in_valid = io_in_valid & _T; // @[ConfigurationMemory.scala 63:44]
  assign neuralNetsweightMatrixMemory_io_in_bits = io_in_bits_wrdata; // @[ConfigurationMemory.scala 61:43]
  assign neuralNetsweightVecMemory_clock = clock;
  assign neuralNetsweightVecMemory_reset = reset;
  assign neuralNetsweightVecMemory_io_in_valid = io_in_valid & _T_2; // @[ConfigurationMemory.scala 75:41]
  assign neuralNetsweightVecMemory_io_in_bits = io_in_bits_wrdata; // @[ConfigurationMemory.scala 73:40]
  assign neuralNetsbiasVecMemory_clock = clock;
  assign neuralNetsbiasVecMemory_reset = reset;
  assign neuralNetsbiasVecMemory_io_in_valid = io_in_valid & _T_4; // @[ConfigurationMemory.scala 86:39]
  assign neuralNetsbiasVecMemory_io_in_bits = io_in_bits_wrdata; // @[ConfigurationMemory.scala 84:38]
  assign neuralNetsbiasScalarMemory_clock = clock;
  assign neuralNetsbiasScalarMemory_reset = reset;
  assign neuralNetsbiasScalarMemory_io_in_valid = io_in_valid & _T_6; // @[ConfigurationMemory.scala 98:42]
  assign neuralNetsbiasScalarMemory_io_in_bits = io_in_bits_wrdata; // @[ConfigurationMemory.scala 96:41]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  inputMuxSel = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      inputMuxSel <= 1'h0;
    end else begin
      if (_T_9) begin
        inputMuxSel <= _T_11;
      end
    end
  end
endmodule
module TLWellnessDataPathBlock(
  input         clock,
  input         reset,
  output        in_ready,
  input         in_valid,
  input  [63:0] in_bits_data,
  input         in_bits_last,
  input         out_ready,
  output        out_valid,
  output [63:0] out_bits_data,
  output        out_bits_last,
  output        in2_ready,
  input         in2_valid,
  input  [63:0] in2_bits_data,
  input         in2_bits_last,
  input         streamIn_valid,
  input  [31:0] streamIn_bits,
  input         streamIn_sync
);
  wire  converter_auto_in_ready; // @[Nodes.scala 106:31]
  wire  converter_auto_in_valid; // @[Nodes.scala 106:31]
  wire [63:0] converter_auto_in_bits_data; // @[Nodes.scala 106:31]
  wire  converter_auto_in_bits_last; // @[Nodes.scala 106:31]
  wire  converter_auto_out_ready; // @[Nodes.scala 106:31]
  wire  converter_auto_out_valid; // @[Nodes.scala 106:31]
  wire [63:0] converter_auto_out_bits_data; // @[Nodes.scala 106:31]
  wire  converter_auto_out_bits_last; // @[Nodes.scala 106:31]
  wire  converter_1_auto_in_ready; // @[Nodes.scala 142:31]
  wire  converter_1_auto_in_valid; // @[Nodes.scala 142:31]
  wire [63:0] converter_1_auto_in_bits_data; // @[Nodes.scala 142:31]
  wire  converter_1_auto_in_bits_last; // @[Nodes.scala 142:31]
  wire  converter_1_auto_out_ready; // @[Nodes.scala 142:31]
  wire  converter_1_auto_out_valid; // @[Nodes.scala 142:31]
  wire [63:0] converter_1_auto_out_bits_data; // @[Nodes.scala 142:31]
  wire  converter_1_auto_out_bits_last; // @[Nodes.scala 142:31]
  wire  converter_2_auto_in_ready; // @[Nodes.scala 142:31]
  wire  converter_2_auto_in_valid; // @[Nodes.scala 142:31]
  wire [63:0] converter_2_auto_in_bits_data; // @[Nodes.scala 142:31]
  wire  converter_2_auto_in_bits_last; // @[Nodes.scala 142:31]
  wire  converter_2_auto_out_ready; // @[Nodes.scala 142:31]
  wire  converter_2_auto_out_valid; // @[Nodes.scala 142:31]
  wire [63:0] converter_2_auto_out_bits_data; // @[Nodes.scala 142:31]
  wire  converter_2_auto_out_bits_last; // @[Nodes.scala 142:31]
  wire  wellness_clock; // @[Wellness.scala 388:26]
  wire  wellness_reset; // @[Wellness.scala 388:26]
  wire  wellness_io_streamIn_valid; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_streamIn_bits; // @[Wellness.scala 388:26]
  wire  wellness_io_in_valid; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_in_bits; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_0_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_0_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_0_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_0_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_1_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_1_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_1_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_1_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_2_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_2_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_2_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_2_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_3_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_3_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_3_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_3_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_4_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_4_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_4_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_4_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_5_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_5_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_5_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_5_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_6_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_6_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_6_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_6_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_7_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_7_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_7_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_7_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_8_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_8_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_8_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_8_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_9_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_9_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_9_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_9_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_10_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_10_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_10_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_10_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_11_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_11_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_11_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_11_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_12_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_12_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_12_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_12_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_13_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_13_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_13_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_13_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_14_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_14_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_14_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_14_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_15_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_15_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_15_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_15_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_16_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_16_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_16_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_16_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_17_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_17_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_17_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_17_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_18_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_18_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_18_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_18_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_19_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_19_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_19_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_19_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_20_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_20_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_20_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_20_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_21_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_21_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_21_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_21_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_22_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_22_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_22_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_22_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_23_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_23_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_23_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_23_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_24_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_24_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_24_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_24_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_25_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_25_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_25_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_25_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_26_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_26_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_26_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_26_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_27_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_27_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_27_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_27_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_28_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_28_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_28_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_28_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_29_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_29_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_29_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_29_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_30_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_30_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_30_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_30_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_31_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_31_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_31_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_31_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_32_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_32_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_32_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_32_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_33_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_33_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_33_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_33_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_34_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_34_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_34_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_34_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_35_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_35_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_35_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_35_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_36_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_36_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_36_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_36_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_37_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_37_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_37_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_37_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_38_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_38_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_38_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_38_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_39_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_39_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_39_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_39_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_40_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_40_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_40_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_40_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_41_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_41_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_41_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_41_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_42_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_42_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_42_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_42_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_43_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_43_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_43_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_43_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_44_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_44_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_44_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_44_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_45_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_45_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_45_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_45_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_46_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_46_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_46_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_46_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_47_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_47_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_47_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_47_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_48_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_48_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_48_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_48_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_49_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_49_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_49_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_49_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_50_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_50_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_50_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_50_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_51_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_51_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_51_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_51_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_52_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_52_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_52_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_52_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_53_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_53_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_53_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_53_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_54_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_54_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_54_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_54_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_55_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_55_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_55_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_55_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_56_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_56_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_56_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_56_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_57_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_57_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_57_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_57_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_58_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_58_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_58_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_58_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_59_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_59_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_59_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_59_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_60_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_60_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_60_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_60_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_61_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_61_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_61_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_61_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_62_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_62_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_62_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_62_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_63_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_63_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_63_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_63_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_64_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_64_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_64_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_64_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_65_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_65_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_65_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_65_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_66_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_66_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_66_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_66_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_67_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_67_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_67_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_67_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_68_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_68_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_68_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_68_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_69_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_69_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_69_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_69_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_70_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_70_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_70_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_70_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_71_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_71_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_71_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_71_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_72_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_72_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_72_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_72_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_73_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_73_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_73_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_73_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_74_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_74_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_74_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_74_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_75_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_75_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_75_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_75_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_76_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_76_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_76_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_76_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_77_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_77_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_77_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_77_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_78_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_78_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_78_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_78_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_79_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_79_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_79_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_79_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_80_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_80_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_80_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_80_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_81_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_81_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_81_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_81_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_82_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_82_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_82_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_82_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_83_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_83_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_83_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_83_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_84_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_84_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_84_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_84_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_85_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_85_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_85_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_85_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_86_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_86_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_86_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_86_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_87_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_87_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_87_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_87_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_88_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_88_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_88_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_88_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_89_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_89_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_89_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_89_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_90_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_90_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_90_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_90_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_91_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_91_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_91_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_91_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_92_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_92_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_92_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_92_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_93_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_93_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_93_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_93_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_94_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_94_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_94_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_94_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_95_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_95_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_95_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_95_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_96_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_96_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_96_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_96_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_97_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_97_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_97_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_97_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_98_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_98_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_98_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_98_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_99_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_99_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_99_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightMatrix_99_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_4; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_5; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_6; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_7; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_8; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_9; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_10; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_11; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_12; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_13; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_14; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_15; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_16; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_17; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_18; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_19; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_20; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_21; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_22; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_23; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_24; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_25; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_26; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_27; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_28; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_29; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_30; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_31; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_32; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_33; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_34; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_35; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_36; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_37; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_38; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_39; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_40; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_41; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_42; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_43; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_44; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_45; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_46; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_47; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_48; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_49; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_50; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_51; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_52; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_53; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_54; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_55; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_56; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_57; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_58; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_59; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_60; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_61; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_62; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_63; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_64; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_65; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_66; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_67; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_68; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_69; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_70; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_71; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_72; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_73; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_74; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_75; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_76; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_77; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_78; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_79; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_80; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_81; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_82; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_83; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_84; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_85; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_86; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_87; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_88; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_89; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_90; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_91; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_92; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_93; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_94; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_95; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_96; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_97; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_98; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsweightVec_99; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_4; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_5; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_6; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_7; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_8; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_9; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_10; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_11; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_12; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_13; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_14; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_15; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_16; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_17; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_18; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_19; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_20; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_21; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_22; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_23; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_24; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_25; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_26; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_27; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_28; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_29; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_30; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_31; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_32; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_33; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_34; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_35; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_36; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_37; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_38; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_39; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_40; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_41; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_42; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_43; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_44; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_45; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_46; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_47; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_48; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_49; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_50; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_51; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_52; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_53; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_54; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_55; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_56; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_57; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_58; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_59; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_60; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_61; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_62; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_63; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_64; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_65; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_66; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_67; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_68; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_69; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_70; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_71; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_72; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_73; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_74; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_75; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_76; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_77; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_78; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_79; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_80; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_81; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_82; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_83; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_84; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_85; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_86; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_87; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_88; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_89; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_90; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_91; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_92; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_93; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_94; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_95; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_96; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_97; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_98; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVec_99; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasScalar_0; // @[Wellness.scala 388:26]
  wire  wellness_io_inConf_bits_confInputMuxSel; // @[Wellness.scala 388:26]
  wire  wellness_io_out_valid; // @[Wellness.scala 388:26]
  wire  wellness_io_out_bits; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_rawVotes; // @[Wellness.scala 388:26]
  wire  configurationMemory_clock; // @[Wellness.scala 398:37]
  wire  configurationMemory_reset; // @[Wellness.scala 398:37]
  wire  configurationMemory_io_in_valid; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_in_bits_wrdata; // @[Wellness.scala 398:37]
  wire [2:0] configurationMemory_io_in_bits_wraddr; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_0_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_0_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_0_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_0_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_1_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_1_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_1_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_1_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_2_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_2_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_2_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_2_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_3_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_3_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_3_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_3_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_4_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_4_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_4_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_4_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_5_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_5_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_5_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_5_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_6_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_6_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_6_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_6_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_7_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_7_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_7_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_7_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_8_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_8_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_8_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_8_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_9_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_9_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_9_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_9_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_10_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_10_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_10_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_10_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_11_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_11_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_11_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_11_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_12_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_12_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_12_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_12_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_13_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_13_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_13_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_13_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_14_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_14_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_14_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_14_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_15_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_15_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_15_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_15_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_16_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_16_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_16_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_16_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_17_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_17_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_17_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_17_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_18_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_18_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_18_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_18_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_19_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_19_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_19_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_19_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_20_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_20_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_20_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_20_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_21_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_21_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_21_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_21_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_22_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_22_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_22_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_22_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_23_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_23_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_23_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_23_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_24_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_24_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_24_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_24_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_25_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_25_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_25_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_25_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_26_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_26_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_26_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_26_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_27_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_27_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_27_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_27_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_28_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_28_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_28_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_28_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_29_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_29_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_29_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_29_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_30_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_30_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_30_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_30_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_31_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_31_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_31_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_31_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_32_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_32_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_32_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_32_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_33_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_33_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_33_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_33_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_34_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_34_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_34_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_34_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_35_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_35_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_35_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_35_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_36_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_36_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_36_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_36_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_37_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_37_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_37_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_37_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_38_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_38_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_38_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_38_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_39_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_39_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_39_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_39_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_40_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_40_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_40_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_40_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_41_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_41_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_41_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_41_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_42_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_42_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_42_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_42_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_43_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_43_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_43_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_43_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_44_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_44_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_44_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_44_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_45_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_45_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_45_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_45_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_46_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_46_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_46_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_46_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_47_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_47_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_47_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_47_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_48_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_48_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_48_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_48_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_49_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_49_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_49_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_49_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_50_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_50_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_50_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_50_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_51_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_51_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_51_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_51_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_52_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_52_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_52_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_52_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_53_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_53_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_53_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_53_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_54_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_54_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_54_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_54_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_55_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_55_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_55_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_55_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_56_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_56_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_56_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_56_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_57_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_57_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_57_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_57_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_58_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_58_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_58_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_58_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_59_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_59_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_59_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_59_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_60_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_60_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_60_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_60_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_61_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_61_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_61_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_61_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_62_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_62_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_62_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_62_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_63_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_63_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_63_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_63_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_64_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_64_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_64_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_64_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_65_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_65_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_65_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_65_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_66_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_66_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_66_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_66_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_67_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_67_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_67_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_67_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_68_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_68_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_68_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_68_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_69_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_69_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_69_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_69_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_70_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_70_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_70_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_70_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_71_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_71_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_71_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_71_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_72_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_72_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_72_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_72_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_73_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_73_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_73_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_73_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_74_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_74_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_74_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_74_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_75_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_75_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_75_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_75_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_76_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_76_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_76_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_76_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_77_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_77_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_77_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_77_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_78_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_78_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_78_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_78_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_79_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_79_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_79_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_79_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_80_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_80_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_80_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_80_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_81_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_81_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_81_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_81_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_82_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_82_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_82_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_82_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_83_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_83_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_83_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_83_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_84_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_84_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_84_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_84_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_85_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_85_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_85_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_85_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_86_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_86_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_86_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_86_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_87_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_87_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_87_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_87_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_88_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_88_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_88_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_88_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_89_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_89_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_89_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_89_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_90_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_90_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_90_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_90_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_91_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_91_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_91_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_91_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_92_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_92_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_92_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_92_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_93_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_93_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_93_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_93_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_94_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_94_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_94_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_94_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_95_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_95_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_95_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_95_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_96_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_96_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_96_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_96_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_97_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_97_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_97_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_97_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_98_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_98_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_98_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_98_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_99_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_99_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_99_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightMatrix_99_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_4; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_5; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_6; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_7; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_8; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_9; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_10; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_11; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_12; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_13; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_14; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_15; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_16; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_17; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_18; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_19; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_20; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_21; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_22; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_23; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_24; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_25; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_26; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_27; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_28; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_29; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_30; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_31; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_32; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_33; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_34; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_35; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_36; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_37; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_38; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_39; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_40; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_41; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_42; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_43; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_44; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_45; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_46; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_47; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_48; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_49; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_50; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_51; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_52; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_53; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_54; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_55; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_56; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_57; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_58; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_59; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_60; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_61; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_62; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_63; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_64; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_65; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_66; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_67; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_68; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_69; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_70; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_71; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_72; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_73; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_74; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_75; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_76; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_77; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_78; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_79; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_80; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_81; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_82; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_83; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_84; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_85; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_86; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_87; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_88; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_89; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_90; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_91; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_92; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_93; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_94; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_95; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_96; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_97; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_98; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsweightVec_99; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_4; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_5; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_6; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_7; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_8; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_9; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_10; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_11; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_12; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_13; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_14; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_15; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_16; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_17; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_18; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_19; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_20; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_21; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_22; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_23; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_24; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_25; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_26; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_27; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_28; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_29; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_30; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_31; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_32; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_33; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_34; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_35; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_36; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_37; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_38; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_39; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_40; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_41; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_42; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_43; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_44; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_45; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_46; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_47; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_48; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_49; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_50; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_51; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_52; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_53; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_54; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_55; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_56; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_57; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_58; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_59; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_60; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_61; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_62; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_63; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_64; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_65; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_66; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_67; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_68; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_69; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_70; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_71; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_72; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_73; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_74; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_75; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_76; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_77; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_78; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_79; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_80; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_81; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_82; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_83; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_84; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_85; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_86; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_87; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_88; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_89; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_90; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_91; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_92; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_93; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_94; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_95; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_96; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_97; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_98; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVec_99; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasScalar_0; // @[Wellness.scala 398:37]
  wire  configurationMemory_io_out_bits_confInputMuxSel; // @[Wellness.scala 398:37]
  wire [63:0] in_1_bits_data; // @[Nodes.scala 333:76 LazyModule.scala 167:31]
  wire [63:0] _T_4; // @[Wellness.scala 408:49]
  wire [31:0] _T_5; // @[Wellness.scala 411:83]
  wire [32:0] _T_6; // @[Cat.scala 30:58]
  wire [63:0] inConf_bits_data; // @[Nodes.scala 333:76 LazyModule.scala 167:31]
  wire [31:0] _T_7; // @[Wellness.scala 418:62]
  wire [31:0] _GEN_0; // @[Wellness.scala 408:49 Wellness.scala 408:49]
  AXI4StreamToBundleBridge converter ( // @[Nodes.scala 106:31]
    .auto_in_ready(converter_auto_in_ready),
    .auto_in_valid(converter_auto_in_valid),
    .auto_in_bits_data(converter_auto_in_bits_data),
    .auto_in_bits_last(converter_auto_in_bits_last),
    .auto_out_ready(converter_auto_out_ready),
    .auto_out_valid(converter_auto_out_valid),
    .auto_out_bits_data(converter_auto_out_bits_data),
    .auto_out_bits_last(converter_auto_out_bits_last)
  );
  AXI4StreamToBundleBridge converter_1 ( // @[Nodes.scala 142:31]
    .auto_in_ready(converter_1_auto_in_ready),
    .auto_in_valid(converter_1_auto_in_valid),
    .auto_in_bits_data(converter_1_auto_in_bits_data),
    .auto_in_bits_last(converter_1_auto_in_bits_last),
    .auto_out_ready(converter_1_auto_out_ready),
    .auto_out_valid(converter_1_auto_out_valid),
    .auto_out_bits_data(converter_1_auto_out_bits_data),
    .auto_out_bits_last(converter_1_auto_out_bits_last)
  );
  AXI4StreamToBundleBridge converter_2 ( // @[Nodes.scala 142:31]
    .auto_in_ready(converter_2_auto_in_ready),
    .auto_in_valid(converter_2_auto_in_valid),
    .auto_in_bits_data(converter_2_auto_in_bits_data),
    .auto_in_bits_last(converter_2_auto_in_bits_last),
    .auto_out_ready(converter_2_auto_out_ready),
    .auto_out_valid(converter_2_auto_out_valid),
    .auto_out_bits_data(converter_2_auto_out_bits_data),
    .auto_out_bits_last(converter_2_auto_out_bits_last)
  );
  WellnessModule wellness ( // @[Wellness.scala 388:26]
    .clock(wellness_clock),
    .reset(wellness_reset),
    .io_streamIn_valid(wellness_io_streamIn_valid),
    .io_streamIn_bits(wellness_io_streamIn_bits),
    .io_in_valid(wellness_io_in_valid),
    .io_in_bits(wellness_io_in_bits),
    .io_inConf_bits_confneuralNetsweightMatrix_0_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_0_0),
    .io_inConf_bits_confneuralNetsweightMatrix_0_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_0_1),
    .io_inConf_bits_confneuralNetsweightMatrix_0_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_0_2),
    .io_inConf_bits_confneuralNetsweightMatrix_0_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_0_3),
    .io_inConf_bits_confneuralNetsweightMatrix_1_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_1_0),
    .io_inConf_bits_confneuralNetsweightMatrix_1_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_1_1),
    .io_inConf_bits_confneuralNetsweightMatrix_1_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_1_2),
    .io_inConf_bits_confneuralNetsweightMatrix_1_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_1_3),
    .io_inConf_bits_confneuralNetsweightMatrix_2_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_2_0),
    .io_inConf_bits_confneuralNetsweightMatrix_2_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_2_1),
    .io_inConf_bits_confneuralNetsweightMatrix_2_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_2_2),
    .io_inConf_bits_confneuralNetsweightMatrix_2_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_2_3),
    .io_inConf_bits_confneuralNetsweightMatrix_3_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_3_0),
    .io_inConf_bits_confneuralNetsweightMatrix_3_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_3_1),
    .io_inConf_bits_confneuralNetsweightMatrix_3_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_3_2),
    .io_inConf_bits_confneuralNetsweightMatrix_3_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_3_3),
    .io_inConf_bits_confneuralNetsweightMatrix_4_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_4_0),
    .io_inConf_bits_confneuralNetsweightMatrix_4_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_4_1),
    .io_inConf_bits_confneuralNetsweightMatrix_4_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_4_2),
    .io_inConf_bits_confneuralNetsweightMatrix_4_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_4_3),
    .io_inConf_bits_confneuralNetsweightMatrix_5_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_5_0),
    .io_inConf_bits_confneuralNetsweightMatrix_5_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_5_1),
    .io_inConf_bits_confneuralNetsweightMatrix_5_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_5_2),
    .io_inConf_bits_confneuralNetsweightMatrix_5_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_5_3),
    .io_inConf_bits_confneuralNetsweightMatrix_6_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_6_0),
    .io_inConf_bits_confneuralNetsweightMatrix_6_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_6_1),
    .io_inConf_bits_confneuralNetsweightMatrix_6_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_6_2),
    .io_inConf_bits_confneuralNetsweightMatrix_6_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_6_3),
    .io_inConf_bits_confneuralNetsweightMatrix_7_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_7_0),
    .io_inConf_bits_confneuralNetsweightMatrix_7_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_7_1),
    .io_inConf_bits_confneuralNetsweightMatrix_7_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_7_2),
    .io_inConf_bits_confneuralNetsweightMatrix_7_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_7_3),
    .io_inConf_bits_confneuralNetsweightMatrix_8_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_8_0),
    .io_inConf_bits_confneuralNetsweightMatrix_8_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_8_1),
    .io_inConf_bits_confneuralNetsweightMatrix_8_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_8_2),
    .io_inConf_bits_confneuralNetsweightMatrix_8_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_8_3),
    .io_inConf_bits_confneuralNetsweightMatrix_9_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_9_0),
    .io_inConf_bits_confneuralNetsweightMatrix_9_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_9_1),
    .io_inConf_bits_confneuralNetsweightMatrix_9_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_9_2),
    .io_inConf_bits_confneuralNetsweightMatrix_9_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_9_3),
    .io_inConf_bits_confneuralNetsweightMatrix_10_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_10_0),
    .io_inConf_bits_confneuralNetsweightMatrix_10_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_10_1),
    .io_inConf_bits_confneuralNetsweightMatrix_10_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_10_2),
    .io_inConf_bits_confneuralNetsweightMatrix_10_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_10_3),
    .io_inConf_bits_confneuralNetsweightMatrix_11_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_11_0),
    .io_inConf_bits_confneuralNetsweightMatrix_11_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_11_1),
    .io_inConf_bits_confneuralNetsweightMatrix_11_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_11_2),
    .io_inConf_bits_confneuralNetsweightMatrix_11_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_11_3),
    .io_inConf_bits_confneuralNetsweightMatrix_12_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_12_0),
    .io_inConf_bits_confneuralNetsweightMatrix_12_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_12_1),
    .io_inConf_bits_confneuralNetsweightMatrix_12_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_12_2),
    .io_inConf_bits_confneuralNetsweightMatrix_12_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_12_3),
    .io_inConf_bits_confneuralNetsweightMatrix_13_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_13_0),
    .io_inConf_bits_confneuralNetsweightMatrix_13_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_13_1),
    .io_inConf_bits_confneuralNetsweightMatrix_13_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_13_2),
    .io_inConf_bits_confneuralNetsweightMatrix_13_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_13_3),
    .io_inConf_bits_confneuralNetsweightMatrix_14_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_14_0),
    .io_inConf_bits_confneuralNetsweightMatrix_14_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_14_1),
    .io_inConf_bits_confneuralNetsweightMatrix_14_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_14_2),
    .io_inConf_bits_confneuralNetsweightMatrix_14_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_14_3),
    .io_inConf_bits_confneuralNetsweightMatrix_15_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_15_0),
    .io_inConf_bits_confneuralNetsweightMatrix_15_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_15_1),
    .io_inConf_bits_confneuralNetsweightMatrix_15_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_15_2),
    .io_inConf_bits_confneuralNetsweightMatrix_15_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_15_3),
    .io_inConf_bits_confneuralNetsweightMatrix_16_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_16_0),
    .io_inConf_bits_confneuralNetsweightMatrix_16_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_16_1),
    .io_inConf_bits_confneuralNetsweightMatrix_16_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_16_2),
    .io_inConf_bits_confneuralNetsweightMatrix_16_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_16_3),
    .io_inConf_bits_confneuralNetsweightMatrix_17_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_17_0),
    .io_inConf_bits_confneuralNetsweightMatrix_17_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_17_1),
    .io_inConf_bits_confneuralNetsweightMatrix_17_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_17_2),
    .io_inConf_bits_confneuralNetsweightMatrix_17_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_17_3),
    .io_inConf_bits_confneuralNetsweightMatrix_18_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_18_0),
    .io_inConf_bits_confneuralNetsweightMatrix_18_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_18_1),
    .io_inConf_bits_confneuralNetsweightMatrix_18_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_18_2),
    .io_inConf_bits_confneuralNetsweightMatrix_18_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_18_3),
    .io_inConf_bits_confneuralNetsweightMatrix_19_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_19_0),
    .io_inConf_bits_confneuralNetsweightMatrix_19_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_19_1),
    .io_inConf_bits_confneuralNetsweightMatrix_19_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_19_2),
    .io_inConf_bits_confneuralNetsweightMatrix_19_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_19_3),
    .io_inConf_bits_confneuralNetsweightMatrix_20_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_20_0),
    .io_inConf_bits_confneuralNetsweightMatrix_20_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_20_1),
    .io_inConf_bits_confneuralNetsweightMatrix_20_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_20_2),
    .io_inConf_bits_confneuralNetsweightMatrix_20_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_20_3),
    .io_inConf_bits_confneuralNetsweightMatrix_21_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_21_0),
    .io_inConf_bits_confneuralNetsweightMatrix_21_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_21_1),
    .io_inConf_bits_confneuralNetsweightMatrix_21_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_21_2),
    .io_inConf_bits_confneuralNetsweightMatrix_21_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_21_3),
    .io_inConf_bits_confneuralNetsweightMatrix_22_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_22_0),
    .io_inConf_bits_confneuralNetsweightMatrix_22_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_22_1),
    .io_inConf_bits_confneuralNetsweightMatrix_22_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_22_2),
    .io_inConf_bits_confneuralNetsweightMatrix_22_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_22_3),
    .io_inConf_bits_confneuralNetsweightMatrix_23_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_23_0),
    .io_inConf_bits_confneuralNetsweightMatrix_23_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_23_1),
    .io_inConf_bits_confneuralNetsweightMatrix_23_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_23_2),
    .io_inConf_bits_confneuralNetsweightMatrix_23_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_23_3),
    .io_inConf_bits_confneuralNetsweightMatrix_24_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_24_0),
    .io_inConf_bits_confneuralNetsweightMatrix_24_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_24_1),
    .io_inConf_bits_confneuralNetsweightMatrix_24_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_24_2),
    .io_inConf_bits_confneuralNetsweightMatrix_24_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_24_3),
    .io_inConf_bits_confneuralNetsweightMatrix_25_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_25_0),
    .io_inConf_bits_confneuralNetsweightMatrix_25_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_25_1),
    .io_inConf_bits_confneuralNetsweightMatrix_25_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_25_2),
    .io_inConf_bits_confneuralNetsweightMatrix_25_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_25_3),
    .io_inConf_bits_confneuralNetsweightMatrix_26_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_26_0),
    .io_inConf_bits_confneuralNetsweightMatrix_26_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_26_1),
    .io_inConf_bits_confneuralNetsweightMatrix_26_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_26_2),
    .io_inConf_bits_confneuralNetsweightMatrix_26_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_26_3),
    .io_inConf_bits_confneuralNetsweightMatrix_27_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_27_0),
    .io_inConf_bits_confneuralNetsweightMatrix_27_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_27_1),
    .io_inConf_bits_confneuralNetsweightMatrix_27_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_27_2),
    .io_inConf_bits_confneuralNetsweightMatrix_27_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_27_3),
    .io_inConf_bits_confneuralNetsweightMatrix_28_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_28_0),
    .io_inConf_bits_confneuralNetsweightMatrix_28_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_28_1),
    .io_inConf_bits_confneuralNetsweightMatrix_28_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_28_2),
    .io_inConf_bits_confneuralNetsweightMatrix_28_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_28_3),
    .io_inConf_bits_confneuralNetsweightMatrix_29_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_29_0),
    .io_inConf_bits_confneuralNetsweightMatrix_29_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_29_1),
    .io_inConf_bits_confneuralNetsweightMatrix_29_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_29_2),
    .io_inConf_bits_confneuralNetsweightMatrix_29_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_29_3),
    .io_inConf_bits_confneuralNetsweightMatrix_30_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_30_0),
    .io_inConf_bits_confneuralNetsweightMatrix_30_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_30_1),
    .io_inConf_bits_confneuralNetsweightMatrix_30_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_30_2),
    .io_inConf_bits_confneuralNetsweightMatrix_30_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_30_3),
    .io_inConf_bits_confneuralNetsweightMatrix_31_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_31_0),
    .io_inConf_bits_confneuralNetsweightMatrix_31_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_31_1),
    .io_inConf_bits_confneuralNetsweightMatrix_31_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_31_2),
    .io_inConf_bits_confneuralNetsweightMatrix_31_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_31_3),
    .io_inConf_bits_confneuralNetsweightMatrix_32_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_32_0),
    .io_inConf_bits_confneuralNetsweightMatrix_32_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_32_1),
    .io_inConf_bits_confneuralNetsweightMatrix_32_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_32_2),
    .io_inConf_bits_confneuralNetsweightMatrix_32_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_32_3),
    .io_inConf_bits_confneuralNetsweightMatrix_33_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_33_0),
    .io_inConf_bits_confneuralNetsweightMatrix_33_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_33_1),
    .io_inConf_bits_confneuralNetsweightMatrix_33_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_33_2),
    .io_inConf_bits_confneuralNetsweightMatrix_33_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_33_3),
    .io_inConf_bits_confneuralNetsweightMatrix_34_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_34_0),
    .io_inConf_bits_confneuralNetsweightMatrix_34_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_34_1),
    .io_inConf_bits_confneuralNetsweightMatrix_34_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_34_2),
    .io_inConf_bits_confneuralNetsweightMatrix_34_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_34_3),
    .io_inConf_bits_confneuralNetsweightMatrix_35_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_35_0),
    .io_inConf_bits_confneuralNetsweightMatrix_35_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_35_1),
    .io_inConf_bits_confneuralNetsweightMatrix_35_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_35_2),
    .io_inConf_bits_confneuralNetsweightMatrix_35_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_35_3),
    .io_inConf_bits_confneuralNetsweightMatrix_36_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_36_0),
    .io_inConf_bits_confneuralNetsweightMatrix_36_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_36_1),
    .io_inConf_bits_confneuralNetsweightMatrix_36_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_36_2),
    .io_inConf_bits_confneuralNetsweightMatrix_36_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_36_3),
    .io_inConf_bits_confneuralNetsweightMatrix_37_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_37_0),
    .io_inConf_bits_confneuralNetsweightMatrix_37_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_37_1),
    .io_inConf_bits_confneuralNetsweightMatrix_37_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_37_2),
    .io_inConf_bits_confneuralNetsweightMatrix_37_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_37_3),
    .io_inConf_bits_confneuralNetsweightMatrix_38_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_38_0),
    .io_inConf_bits_confneuralNetsweightMatrix_38_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_38_1),
    .io_inConf_bits_confneuralNetsweightMatrix_38_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_38_2),
    .io_inConf_bits_confneuralNetsweightMatrix_38_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_38_3),
    .io_inConf_bits_confneuralNetsweightMatrix_39_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_39_0),
    .io_inConf_bits_confneuralNetsweightMatrix_39_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_39_1),
    .io_inConf_bits_confneuralNetsweightMatrix_39_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_39_2),
    .io_inConf_bits_confneuralNetsweightMatrix_39_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_39_3),
    .io_inConf_bits_confneuralNetsweightMatrix_40_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_40_0),
    .io_inConf_bits_confneuralNetsweightMatrix_40_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_40_1),
    .io_inConf_bits_confneuralNetsweightMatrix_40_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_40_2),
    .io_inConf_bits_confneuralNetsweightMatrix_40_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_40_3),
    .io_inConf_bits_confneuralNetsweightMatrix_41_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_41_0),
    .io_inConf_bits_confneuralNetsweightMatrix_41_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_41_1),
    .io_inConf_bits_confneuralNetsweightMatrix_41_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_41_2),
    .io_inConf_bits_confneuralNetsweightMatrix_41_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_41_3),
    .io_inConf_bits_confneuralNetsweightMatrix_42_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_42_0),
    .io_inConf_bits_confneuralNetsweightMatrix_42_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_42_1),
    .io_inConf_bits_confneuralNetsweightMatrix_42_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_42_2),
    .io_inConf_bits_confneuralNetsweightMatrix_42_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_42_3),
    .io_inConf_bits_confneuralNetsweightMatrix_43_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_43_0),
    .io_inConf_bits_confneuralNetsweightMatrix_43_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_43_1),
    .io_inConf_bits_confneuralNetsweightMatrix_43_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_43_2),
    .io_inConf_bits_confneuralNetsweightMatrix_43_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_43_3),
    .io_inConf_bits_confneuralNetsweightMatrix_44_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_44_0),
    .io_inConf_bits_confneuralNetsweightMatrix_44_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_44_1),
    .io_inConf_bits_confneuralNetsweightMatrix_44_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_44_2),
    .io_inConf_bits_confneuralNetsweightMatrix_44_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_44_3),
    .io_inConf_bits_confneuralNetsweightMatrix_45_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_45_0),
    .io_inConf_bits_confneuralNetsweightMatrix_45_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_45_1),
    .io_inConf_bits_confneuralNetsweightMatrix_45_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_45_2),
    .io_inConf_bits_confneuralNetsweightMatrix_45_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_45_3),
    .io_inConf_bits_confneuralNetsweightMatrix_46_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_46_0),
    .io_inConf_bits_confneuralNetsweightMatrix_46_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_46_1),
    .io_inConf_bits_confneuralNetsweightMatrix_46_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_46_2),
    .io_inConf_bits_confneuralNetsweightMatrix_46_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_46_3),
    .io_inConf_bits_confneuralNetsweightMatrix_47_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_47_0),
    .io_inConf_bits_confneuralNetsweightMatrix_47_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_47_1),
    .io_inConf_bits_confneuralNetsweightMatrix_47_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_47_2),
    .io_inConf_bits_confneuralNetsweightMatrix_47_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_47_3),
    .io_inConf_bits_confneuralNetsweightMatrix_48_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_48_0),
    .io_inConf_bits_confneuralNetsweightMatrix_48_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_48_1),
    .io_inConf_bits_confneuralNetsweightMatrix_48_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_48_2),
    .io_inConf_bits_confneuralNetsweightMatrix_48_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_48_3),
    .io_inConf_bits_confneuralNetsweightMatrix_49_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_49_0),
    .io_inConf_bits_confneuralNetsweightMatrix_49_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_49_1),
    .io_inConf_bits_confneuralNetsweightMatrix_49_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_49_2),
    .io_inConf_bits_confneuralNetsweightMatrix_49_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_49_3),
    .io_inConf_bits_confneuralNetsweightMatrix_50_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_50_0),
    .io_inConf_bits_confneuralNetsweightMatrix_50_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_50_1),
    .io_inConf_bits_confneuralNetsweightMatrix_50_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_50_2),
    .io_inConf_bits_confneuralNetsweightMatrix_50_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_50_3),
    .io_inConf_bits_confneuralNetsweightMatrix_51_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_51_0),
    .io_inConf_bits_confneuralNetsweightMatrix_51_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_51_1),
    .io_inConf_bits_confneuralNetsweightMatrix_51_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_51_2),
    .io_inConf_bits_confneuralNetsweightMatrix_51_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_51_3),
    .io_inConf_bits_confneuralNetsweightMatrix_52_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_52_0),
    .io_inConf_bits_confneuralNetsweightMatrix_52_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_52_1),
    .io_inConf_bits_confneuralNetsweightMatrix_52_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_52_2),
    .io_inConf_bits_confneuralNetsweightMatrix_52_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_52_3),
    .io_inConf_bits_confneuralNetsweightMatrix_53_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_53_0),
    .io_inConf_bits_confneuralNetsweightMatrix_53_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_53_1),
    .io_inConf_bits_confneuralNetsweightMatrix_53_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_53_2),
    .io_inConf_bits_confneuralNetsweightMatrix_53_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_53_3),
    .io_inConf_bits_confneuralNetsweightMatrix_54_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_54_0),
    .io_inConf_bits_confneuralNetsweightMatrix_54_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_54_1),
    .io_inConf_bits_confneuralNetsweightMatrix_54_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_54_2),
    .io_inConf_bits_confneuralNetsweightMatrix_54_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_54_3),
    .io_inConf_bits_confneuralNetsweightMatrix_55_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_55_0),
    .io_inConf_bits_confneuralNetsweightMatrix_55_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_55_1),
    .io_inConf_bits_confneuralNetsweightMatrix_55_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_55_2),
    .io_inConf_bits_confneuralNetsweightMatrix_55_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_55_3),
    .io_inConf_bits_confneuralNetsweightMatrix_56_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_56_0),
    .io_inConf_bits_confneuralNetsweightMatrix_56_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_56_1),
    .io_inConf_bits_confneuralNetsweightMatrix_56_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_56_2),
    .io_inConf_bits_confneuralNetsweightMatrix_56_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_56_3),
    .io_inConf_bits_confneuralNetsweightMatrix_57_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_57_0),
    .io_inConf_bits_confneuralNetsweightMatrix_57_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_57_1),
    .io_inConf_bits_confneuralNetsweightMatrix_57_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_57_2),
    .io_inConf_bits_confneuralNetsweightMatrix_57_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_57_3),
    .io_inConf_bits_confneuralNetsweightMatrix_58_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_58_0),
    .io_inConf_bits_confneuralNetsweightMatrix_58_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_58_1),
    .io_inConf_bits_confneuralNetsweightMatrix_58_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_58_2),
    .io_inConf_bits_confneuralNetsweightMatrix_58_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_58_3),
    .io_inConf_bits_confneuralNetsweightMatrix_59_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_59_0),
    .io_inConf_bits_confneuralNetsweightMatrix_59_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_59_1),
    .io_inConf_bits_confneuralNetsweightMatrix_59_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_59_2),
    .io_inConf_bits_confneuralNetsweightMatrix_59_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_59_3),
    .io_inConf_bits_confneuralNetsweightMatrix_60_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_60_0),
    .io_inConf_bits_confneuralNetsweightMatrix_60_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_60_1),
    .io_inConf_bits_confneuralNetsweightMatrix_60_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_60_2),
    .io_inConf_bits_confneuralNetsweightMatrix_60_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_60_3),
    .io_inConf_bits_confneuralNetsweightMatrix_61_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_61_0),
    .io_inConf_bits_confneuralNetsweightMatrix_61_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_61_1),
    .io_inConf_bits_confneuralNetsweightMatrix_61_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_61_2),
    .io_inConf_bits_confneuralNetsweightMatrix_61_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_61_3),
    .io_inConf_bits_confneuralNetsweightMatrix_62_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_62_0),
    .io_inConf_bits_confneuralNetsweightMatrix_62_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_62_1),
    .io_inConf_bits_confneuralNetsweightMatrix_62_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_62_2),
    .io_inConf_bits_confneuralNetsweightMatrix_62_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_62_3),
    .io_inConf_bits_confneuralNetsweightMatrix_63_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_63_0),
    .io_inConf_bits_confneuralNetsweightMatrix_63_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_63_1),
    .io_inConf_bits_confneuralNetsweightMatrix_63_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_63_2),
    .io_inConf_bits_confneuralNetsweightMatrix_63_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_63_3),
    .io_inConf_bits_confneuralNetsweightMatrix_64_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_64_0),
    .io_inConf_bits_confneuralNetsweightMatrix_64_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_64_1),
    .io_inConf_bits_confneuralNetsweightMatrix_64_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_64_2),
    .io_inConf_bits_confneuralNetsweightMatrix_64_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_64_3),
    .io_inConf_bits_confneuralNetsweightMatrix_65_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_65_0),
    .io_inConf_bits_confneuralNetsweightMatrix_65_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_65_1),
    .io_inConf_bits_confneuralNetsweightMatrix_65_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_65_2),
    .io_inConf_bits_confneuralNetsweightMatrix_65_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_65_3),
    .io_inConf_bits_confneuralNetsweightMatrix_66_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_66_0),
    .io_inConf_bits_confneuralNetsweightMatrix_66_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_66_1),
    .io_inConf_bits_confneuralNetsweightMatrix_66_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_66_2),
    .io_inConf_bits_confneuralNetsweightMatrix_66_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_66_3),
    .io_inConf_bits_confneuralNetsweightMatrix_67_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_67_0),
    .io_inConf_bits_confneuralNetsweightMatrix_67_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_67_1),
    .io_inConf_bits_confneuralNetsweightMatrix_67_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_67_2),
    .io_inConf_bits_confneuralNetsweightMatrix_67_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_67_3),
    .io_inConf_bits_confneuralNetsweightMatrix_68_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_68_0),
    .io_inConf_bits_confneuralNetsweightMatrix_68_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_68_1),
    .io_inConf_bits_confneuralNetsweightMatrix_68_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_68_2),
    .io_inConf_bits_confneuralNetsweightMatrix_68_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_68_3),
    .io_inConf_bits_confneuralNetsweightMatrix_69_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_69_0),
    .io_inConf_bits_confneuralNetsweightMatrix_69_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_69_1),
    .io_inConf_bits_confneuralNetsweightMatrix_69_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_69_2),
    .io_inConf_bits_confneuralNetsweightMatrix_69_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_69_3),
    .io_inConf_bits_confneuralNetsweightMatrix_70_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_70_0),
    .io_inConf_bits_confneuralNetsweightMatrix_70_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_70_1),
    .io_inConf_bits_confneuralNetsweightMatrix_70_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_70_2),
    .io_inConf_bits_confneuralNetsweightMatrix_70_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_70_3),
    .io_inConf_bits_confneuralNetsweightMatrix_71_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_71_0),
    .io_inConf_bits_confneuralNetsweightMatrix_71_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_71_1),
    .io_inConf_bits_confneuralNetsweightMatrix_71_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_71_2),
    .io_inConf_bits_confneuralNetsweightMatrix_71_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_71_3),
    .io_inConf_bits_confneuralNetsweightMatrix_72_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_72_0),
    .io_inConf_bits_confneuralNetsweightMatrix_72_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_72_1),
    .io_inConf_bits_confneuralNetsweightMatrix_72_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_72_2),
    .io_inConf_bits_confneuralNetsweightMatrix_72_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_72_3),
    .io_inConf_bits_confneuralNetsweightMatrix_73_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_73_0),
    .io_inConf_bits_confneuralNetsweightMatrix_73_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_73_1),
    .io_inConf_bits_confneuralNetsweightMatrix_73_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_73_2),
    .io_inConf_bits_confneuralNetsweightMatrix_73_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_73_3),
    .io_inConf_bits_confneuralNetsweightMatrix_74_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_74_0),
    .io_inConf_bits_confneuralNetsweightMatrix_74_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_74_1),
    .io_inConf_bits_confneuralNetsweightMatrix_74_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_74_2),
    .io_inConf_bits_confneuralNetsweightMatrix_74_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_74_3),
    .io_inConf_bits_confneuralNetsweightMatrix_75_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_75_0),
    .io_inConf_bits_confneuralNetsweightMatrix_75_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_75_1),
    .io_inConf_bits_confneuralNetsweightMatrix_75_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_75_2),
    .io_inConf_bits_confneuralNetsweightMatrix_75_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_75_3),
    .io_inConf_bits_confneuralNetsweightMatrix_76_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_76_0),
    .io_inConf_bits_confneuralNetsweightMatrix_76_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_76_1),
    .io_inConf_bits_confneuralNetsweightMatrix_76_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_76_2),
    .io_inConf_bits_confneuralNetsweightMatrix_76_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_76_3),
    .io_inConf_bits_confneuralNetsweightMatrix_77_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_77_0),
    .io_inConf_bits_confneuralNetsweightMatrix_77_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_77_1),
    .io_inConf_bits_confneuralNetsweightMatrix_77_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_77_2),
    .io_inConf_bits_confneuralNetsweightMatrix_77_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_77_3),
    .io_inConf_bits_confneuralNetsweightMatrix_78_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_78_0),
    .io_inConf_bits_confneuralNetsweightMatrix_78_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_78_1),
    .io_inConf_bits_confneuralNetsweightMatrix_78_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_78_2),
    .io_inConf_bits_confneuralNetsweightMatrix_78_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_78_3),
    .io_inConf_bits_confneuralNetsweightMatrix_79_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_79_0),
    .io_inConf_bits_confneuralNetsweightMatrix_79_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_79_1),
    .io_inConf_bits_confneuralNetsweightMatrix_79_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_79_2),
    .io_inConf_bits_confneuralNetsweightMatrix_79_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_79_3),
    .io_inConf_bits_confneuralNetsweightMatrix_80_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_80_0),
    .io_inConf_bits_confneuralNetsweightMatrix_80_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_80_1),
    .io_inConf_bits_confneuralNetsweightMatrix_80_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_80_2),
    .io_inConf_bits_confneuralNetsweightMatrix_80_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_80_3),
    .io_inConf_bits_confneuralNetsweightMatrix_81_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_81_0),
    .io_inConf_bits_confneuralNetsweightMatrix_81_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_81_1),
    .io_inConf_bits_confneuralNetsweightMatrix_81_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_81_2),
    .io_inConf_bits_confneuralNetsweightMatrix_81_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_81_3),
    .io_inConf_bits_confneuralNetsweightMatrix_82_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_82_0),
    .io_inConf_bits_confneuralNetsweightMatrix_82_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_82_1),
    .io_inConf_bits_confneuralNetsweightMatrix_82_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_82_2),
    .io_inConf_bits_confneuralNetsweightMatrix_82_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_82_3),
    .io_inConf_bits_confneuralNetsweightMatrix_83_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_83_0),
    .io_inConf_bits_confneuralNetsweightMatrix_83_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_83_1),
    .io_inConf_bits_confneuralNetsweightMatrix_83_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_83_2),
    .io_inConf_bits_confneuralNetsweightMatrix_83_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_83_3),
    .io_inConf_bits_confneuralNetsweightMatrix_84_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_84_0),
    .io_inConf_bits_confneuralNetsweightMatrix_84_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_84_1),
    .io_inConf_bits_confneuralNetsweightMatrix_84_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_84_2),
    .io_inConf_bits_confneuralNetsweightMatrix_84_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_84_3),
    .io_inConf_bits_confneuralNetsweightMatrix_85_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_85_0),
    .io_inConf_bits_confneuralNetsweightMatrix_85_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_85_1),
    .io_inConf_bits_confneuralNetsweightMatrix_85_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_85_2),
    .io_inConf_bits_confneuralNetsweightMatrix_85_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_85_3),
    .io_inConf_bits_confneuralNetsweightMatrix_86_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_86_0),
    .io_inConf_bits_confneuralNetsweightMatrix_86_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_86_1),
    .io_inConf_bits_confneuralNetsweightMatrix_86_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_86_2),
    .io_inConf_bits_confneuralNetsweightMatrix_86_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_86_3),
    .io_inConf_bits_confneuralNetsweightMatrix_87_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_87_0),
    .io_inConf_bits_confneuralNetsweightMatrix_87_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_87_1),
    .io_inConf_bits_confneuralNetsweightMatrix_87_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_87_2),
    .io_inConf_bits_confneuralNetsweightMatrix_87_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_87_3),
    .io_inConf_bits_confneuralNetsweightMatrix_88_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_88_0),
    .io_inConf_bits_confneuralNetsweightMatrix_88_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_88_1),
    .io_inConf_bits_confneuralNetsweightMatrix_88_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_88_2),
    .io_inConf_bits_confneuralNetsweightMatrix_88_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_88_3),
    .io_inConf_bits_confneuralNetsweightMatrix_89_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_89_0),
    .io_inConf_bits_confneuralNetsweightMatrix_89_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_89_1),
    .io_inConf_bits_confneuralNetsweightMatrix_89_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_89_2),
    .io_inConf_bits_confneuralNetsweightMatrix_89_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_89_3),
    .io_inConf_bits_confneuralNetsweightMatrix_90_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_90_0),
    .io_inConf_bits_confneuralNetsweightMatrix_90_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_90_1),
    .io_inConf_bits_confneuralNetsweightMatrix_90_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_90_2),
    .io_inConf_bits_confneuralNetsweightMatrix_90_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_90_3),
    .io_inConf_bits_confneuralNetsweightMatrix_91_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_91_0),
    .io_inConf_bits_confneuralNetsweightMatrix_91_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_91_1),
    .io_inConf_bits_confneuralNetsweightMatrix_91_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_91_2),
    .io_inConf_bits_confneuralNetsweightMatrix_91_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_91_3),
    .io_inConf_bits_confneuralNetsweightMatrix_92_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_92_0),
    .io_inConf_bits_confneuralNetsweightMatrix_92_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_92_1),
    .io_inConf_bits_confneuralNetsweightMatrix_92_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_92_2),
    .io_inConf_bits_confneuralNetsweightMatrix_92_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_92_3),
    .io_inConf_bits_confneuralNetsweightMatrix_93_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_93_0),
    .io_inConf_bits_confneuralNetsweightMatrix_93_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_93_1),
    .io_inConf_bits_confneuralNetsweightMatrix_93_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_93_2),
    .io_inConf_bits_confneuralNetsweightMatrix_93_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_93_3),
    .io_inConf_bits_confneuralNetsweightMatrix_94_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_94_0),
    .io_inConf_bits_confneuralNetsweightMatrix_94_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_94_1),
    .io_inConf_bits_confneuralNetsweightMatrix_94_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_94_2),
    .io_inConf_bits_confneuralNetsweightMatrix_94_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_94_3),
    .io_inConf_bits_confneuralNetsweightMatrix_95_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_95_0),
    .io_inConf_bits_confneuralNetsweightMatrix_95_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_95_1),
    .io_inConf_bits_confneuralNetsweightMatrix_95_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_95_2),
    .io_inConf_bits_confneuralNetsweightMatrix_95_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_95_3),
    .io_inConf_bits_confneuralNetsweightMatrix_96_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_96_0),
    .io_inConf_bits_confneuralNetsweightMatrix_96_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_96_1),
    .io_inConf_bits_confneuralNetsweightMatrix_96_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_96_2),
    .io_inConf_bits_confneuralNetsweightMatrix_96_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_96_3),
    .io_inConf_bits_confneuralNetsweightMatrix_97_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_97_0),
    .io_inConf_bits_confneuralNetsweightMatrix_97_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_97_1),
    .io_inConf_bits_confneuralNetsweightMatrix_97_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_97_2),
    .io_inConf_bits_confneuralNetsweightMatrix_97_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_97_3),
    .io_inConf_bits_confneuralNetsweightMatrix_98_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_98_0),
    .io_inConf_bits_confneuralNetsweightMatrix_98_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_98_1),
    .io_inConf_bits_confneuralNetsweightMatrix_98_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_98_2),
    .io_inConf_bits_confneuralNetsweightMatrix_98_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_98_3),
    .io_inConf_bits_confneuralNetsweightMatrix_99_0(wellness_io_inConf_bits_confneuralNetsweightMatrix_99_0),
    .io_inConf_bits_confneuralNetsweightMatrix_99_1(wellness_io_inConf_bits_confneuralNetsweightMatrix_99_1),
    .io_inConf_bits_confneuralNetsweightMatrix_99_2(wellness_io_inConf_bits_confneuralNetsweightMatrix_99_2),
    .io_inConf_bits_confneuralNetsweightMatrix_99_3(wellness_io_inConf_bits_confneuralNetsweightMatrix_99_3),
    .io_inConf_bits_confneuralNetsweightVec_0(wellness_io_inConf_bits_confneuralNetsweightVec_0),
    .io_inConf_bits_confneuralNetsweightVec_1(wellness_io_inConf_bits_confneuralNetsweightVec_1),
    .io_inConf_bits_confneuralNetsweightVec_2(wellness_io_inConf_bits_confneuralNetsweightVec_2),
    .io_inConf_bits_confneuralNetsweightVec_3(wellness_io_inConf_bits_confneuralNetsweightVec_3),
    .io_inConf_bits_confneuralNetsweightVec_4(wellness_io_inConf_bits_confneuralNetsweightVec_4),
    .io_inConf_bits_confneuralNetsweightVec_5(wellness_io_inConf_bits_confneuralNetsweightVec_5),
    .io_inConf_bits_confneuralNetsweightVec_6(wellness_io_inConf_bits_confneuralNetsweightVec_6),
    .io_inConf_bits_confneuralNetsweightVec_7(wellness_io_inConf_bits_confneuralNetsweightVec_7),
    .io_inConf_bits_confneuralNetsweightVec_8(wellness_io_inConf_bits_confneuralNetsweightVec_8),
    .io_inConf_bits_confneuralNetsweightVec_9(wellness_io_inConf_bits_confneuralNetsweightVec_9),
    .io_inConf_bits_confneuralNetsweightVec_10(wellness_io_inConf_bits_confneuralNetsweightVec_10),
    .io_inConf_bits_confneuralNetsweightVec_11(wellness_io_inConf_bits_confneuralNetsweightVec_11),
    .io_inConf_bits_confneuralNetsweightVec_12(wellness_io_inConf_bits_confneuralNetsweightVec_12),
    .io_inConf_bits_confneuralNetsweightVec_13(wellness_io_inConf_bits_confneuralNetsweightVec_13),
    .io_inConf_bits_confneuralNetsweightVec_14(wellness_io_inConf_bits_confneuralNetsweightVec_14),
    .io_inConf_bits_confneuralNetsweightVec_15(wellness_io_inConf_bits_confneuralNetsweightVec_15),
    .io_inConf_bits_confneuralNetsweightVec_16(wellness_io_inConf_bits_confneuralNetsweightVec_16),
    .io_inConf_bits_confneuralNetsweightVec_17(wellness_io_inConf_bits_confneuralNetsweightVec_17),
    .io_inConf_bits_confneuralNetsweightVec_18(wellness_io_inConf_bits_confneuralNetsweightVec_18),
    .io_inConf_bits_confneuralNetsweightVec_19(wellness_io_inConf_bits_confneuralNetsweightVec_19),
    .io_inConf_bits_confneuralNetsweightVec_20(wellness_io_inConf_bits_confneuralNetsweightVec_20),
    .io_inConf_bits_confneuralNetsweightVec_21(wellness_io_inConf_bits_confneuralNetsweightVec_21),
    .io_inConf_bits_confneuralNetsweightVec_22(wellness_io_inConf_bits_confneuralNetsweightVec_22),
    .io_inConf_bits_confneuralNetsweightVec_23(wellness_io_inConf_bits_confneuralNetsweightVec_23),
    .io_inConf_bits_confneuralNetsweightVec_24(wellness_io_inConf_bits_confneuralNetsweightVec_24),
    .io_inConf_bits_confneuralNetsweightVec_25(wellness_io_inConf_bits_confneuralNetsweightVec_25),
    .io_inConf_bits_confneuralNetsweightVec_26(wellness_io_inConf_bits_confneuralNetsweightVec_26),
    .io_inConf_bits_confneuralNetsweightVec_27(wellness_io_inConf_bits_confneuralNetsweightVec_27),
    .io_inConf_bits_confneuralNetsweightVec_28(wellness_io_inConf_bits_confneuralNetsweightVec_28),
    .io_inConf_bits_confneuralNetsweightVec_29(wellness_io_inConf_bits_confneuralNetsweightVec_29),
    .io_inConf_bits_confneuralNetsweightVec_30(wellness_io_inConf_bits_confneuralNetsweightVec_30),
    .io_inConf_bits_confneuralNetsweightVec_31(wellness_io_inConf_bits_confneuralNetsweightVec_31),
    .io_inConf_bits_confneuralNetsweightVec_32(wellness_io_inConf_bits_confneuralNetsweightVec_32),
    .io_inConf_bits_confneuralNetsweightVec_33(wellness_io_inConf_bits_confneuralNetsweightVec_33),
    .io_inConf_bits_confneuralNetsweightVec_34(wellness_io_inConf_bits_confneuralNetsweightVec_34),
    .io_inConf_bits_confneuralNetsweightVec_35(wellness_io_inConf_bits_confneuralNetsweightVec_35),
    .io_inConf_bits_confneuralNetsweightVec_36(wellness_io_inConf_bits_confneuralNetsweightVec_36),
    .io_inConf_bits_confneuralNetsweightVec_37(wellness_io_inConf_bits_confneuralNetsweightVec_37),
    .io_inConf_bits_confneuralNetsweightVec_38(wellness_io_inConf_bits_confneuralNetsweightVec_38),
    .io_inConf_bits_confneuralNetsweightVec_39(wellness_io_inConf_bits_confneuralNetsweightVec_39),
    .io_inConf_bits_confneuralNetsweightVec_40(wellness_io_inConf_bits_confneuralNetsweightVec_40),
    .io_inConf_bits_confneuralNetsweightVec_41(wellness_io_inConf_bits_confneuralNetsweightVec_41),
    .io_inConf_bits_confneuralNetsweightVec_42(wellness_io_inConf_bits_confneuralNetsweightVec_42),
    .io_inConf_bits_confneuralNetsweightVec_43(wellness_io_inConf_bits_confneuralNetsweightVec_43),
    .io_inConf_bits_confneuralNetsweightVec_44(wellness_io_inConf_bits_confneuralNetsweightVec_44),
    .io_inConf_bits_confneuralNetsweightVec_45(wellness_io_inConf_bits_confneuralNetsweightVec_45),
    .io_inConf_bits_confneuralNetsweightVec_46(wellness_io_inConf_bits_confneuralNetsweightVec_46),
    .io_inConf_bits_confneuralNetsweightVec_47(wellness_io_inConf_bits_confneuralNetsweightVec_47),
    .io_inConf_bits_confneuralNetsweightVec_48(wellness_io_inConf_bits_confneuralNetsweightVec_48),
    .io_inConf_bits_confneuralNetsweightVec_49(wellness_io_inConf_bits_confneuralNetsweightVec_49),
    .io_inConf_bits_confneuralNetsweightVec_50(wellness_io_inConf_bits_confneuralNetsweightVec_50),
    .io_inConf_bits_confneuralNetsweightVec_51(wellness_io_inConf_bits_confneuralNetsweightVec_51),
    .io_inConf_bits_confneuralNetsweightVec_52(wellness_io_inConf_bits_confneuralNetsweightVec_52),
    .io_inConf_bits_confneuralNetsweightVec_53(wellness_io_inConf_bits_confneuralNetsweightVec_53),
    .io_inConf_bits_confneuralNetsweightVec_54(wellness_io_inConf_bits_confneuralNetsweightVec_54),
    .io_inConf_bits_confneuralNetsweightVec_55(wellness_io_inConf_bits_confneuralNetsweightVec_55),
    .io_inConf_bits_confneuralNetsweightVec_56(wellness_io_inConf_bits_confneuralNetsweightVec_56),
    .io_inConf_bits_confneuralNetsweightVec_57(wellness_io_inConf_bits_confneuralNetsweightVec_57),
    .io_inConf_bits_confneuralNetsweightVec_58(wellness_io_inConf_bits_confneuralNetsweightVec_58),
    .io_inConf_bits_confneuralNetsweightVec_59(wellness_io_inConf_bits_confneuralNetsweightVec_59),
    .io_inConf_bits_confneuralNetsweightVec_60(wellness_io_inConf_bits_confneuralNetsweightVec_60),
    .io_inConf_bits_confneuralNetsweightVec_61(wellness_io_inConf_bits_confneuralNetsweightVec_61),
    .io_inConf_bits_confneuralNetsweightVec_62(wellness_io_inConf_bits_confneuralNetsweightVec_62),
    .io_inConf_bits_confneuralNetsweightVec_63(wellness_io_inConf_bits_confneuralNetsweightVec_63),
    .io_inConf_bits_confneuralNetsweightVec_64(wellness_io_inConf_bits_confneuralNetsweightVec_64),
    .io_inConf_bits_confneuralNetsweightVec_65(wellness_io_inConf_bits_confneuralNetsweightVec_65),
    .io_inConf_bits_confneuralNetsweightVec_66(wellness_io_inConf_bits_confneuralNetsweightVec_66),
    .io_inConf_bits_confneuralNetsweightVec_67(wellness_io_inConf_bits_confneuralNetsweightVec_67),
    .io_inConf_bits_confneuralNetsweightVec_68(wellness_io_inConf_bits_confneuralNetsweightVec_68),
    .io_inConf_bits_confneuralNetsweightVec_69(wellness_io_inConf_bits_confneuralNetsweightVec_69),
    .io_inConf_bits_confneuralNetsweightVec_70(wellness_io_inConf_bits_confneuralNetsweightVec_70),
    .io_inConf_bits_confneuralNetsweightVec_71(wellness_io_inConf_bits_confneuralNetsweightVec_71),
    .io_inConf_bits_confneuralNetsweightVec_72(wellness_io_inConf_bits_confneuralNetsweightVec_72),
    .io_inConf_bits_confneuralNetsweightVec_73(wellness_io_inConf_bits_confneuralNetsweightVec_73),
    .io_inConf_bits_confneuralNetsweightVec_74(wellness_io_inConf_bits_confneuralNetsweightVec_74),
    .io_inConf_bits_confneuralNetsweightVec_75(wellness_io_inConf_bits_confneuralNetsweightVec_75),
    .io_inConf_bits_confneuralNetsweightVec_76(wellness_io_inConf_bits_confneuralNetsweightVec_76),
    .io_inConf_bits_confneuralNetsweightVec_77(wellness_io_inConf_bits_confneuralNetsweightVec_77),
    .io_inConf_bits_confneuralNetsweightVec_78(wellness_io_inConf_bits_confneuralNetsweightVec_78),
    .io_inConf_bits_confneuralNetsweightVec_79(wellness_io_inConf_bits_confneuralNetsweightVec_79),
    .io_inConf_bits_confneuralNetsweightVec_80(wellness_io_inConf_bits_confneuralNetsweightVec_80),
    .io_inConf_bits_confneuralNetsweightVec_81(wellness_io_inConf_bits_confneuralNetsweightVec_81),
    .io_inConf_bits_confneuralNetsweightVec_82(wellness_io_inConf_bits_confneuralNetsweightVec_82),
    .io_inConf_bits_confneuralNetsweightVec_83(wellness_io_inConf_bits_confneuralNetsweightVec_83),
    .io_inConf_bits_confneuralNetsweightVec_84(wellness_io_inConf_bits_confneuralNetsweightVec_84),
    .io_inConf_bits_confneuralNetsweightVec_85(wellness_io_inConf_bits_confneuralNetsweightVec_85),
    .io_inConf_bits_confneuralNetsweightVec_86(wellness_io_inConf_bits_confneuralNetsweightVec_86),
    .io_inConf_bits_confneuralNetsweightVec_87(wellness_io_inConf_bits_confneuralNetsweightVec_87),
    .io_inConf_bits_confneuralNetsweightVec_88(wellness_io_inConf_bits_confneuralNetsweightVec_88),
    .io_inConf_bits_confneuralNetsweightVec_89(wellness_io_inConf_bits_confneuralNetsweightVec_89),
    .io_inConf_bits_confneuralNetsweightVec_90(wellness_io_inConf_bits_confneuralNetsweightVec_90),
    .io_inConf_bits_confneuralNetsweightVec_91(wellness_io_inConf_bits_confneuralNetsweightVec_91),
    .io_inConf_bits_confneuralNetsweightVec_92(wellness_io_inConf_bits_confneuralNetsweightVec_92),
    .io_inConf_bits_confneuralNetsweightVec_93(wellness_io_inConf_bits_confneuralNetsweightVec_93),
    .io_inConf_bits_confneuralNetsweightVec_94(wellness_io_inConf_bits_confneuralNetsweightVec_94),
    .io_inConf_bits_confneuralNetsweightVec_95(wellness_io_inConf_bits_confneuralNetsweightVec_95),
    .io_inConf_bits_confneuralNetsweightVec_96(wellness_io_inConf_bits_confneuralNetsweightVec_96),
    .io_inConf_bits_confneuralNetsweightVec_97(wellness_io_inConf_bits_confneuralNetsweightVec_97),
    .io_inConf_bits_confneuralNetsweightVec_98(wellness_io_inConf_bits_confneuralNetsweightVec_98),
    .io_inConf_bits_confneuralNetsweightVec_99(wellness_io_inConf_bits_confneuralNetsweightVec_99),
    .io_inConf_bits_confneuralNetsbiasVec_0(wellness_io_inConf_bits_confneuralNetsbiasVec_0),
    .io_inConf_bits_confneuralNetsbiasVec_1(wellness_io_inConf_bits_confneuralNetsbiasVec_1),
    .io_inConf_bits_confneuralNetsbiasVec_2(wellness_io_inConf_bits_confneuralNetsbiasVec_2),
    .io_inConf_bits_confneuralNetsbiasVec_3(wellness_io_inConf_bits_confneuralNetsbiasVec_3),
    .io_inConf_bits_confneuralNetsbiasVec_4(wellness_io_inConf_bits_confneuralNetsbiasVec_4),
    .io_inConf_bits_confneuralNetsbiasVec_5(wellness_io_inConf_bits_confneuralNetsbiasVec_5),
    .io_inConf_bits_confneuralNetsbiasVec_6(wellness_io_inConf_bits_confneuralNetsbiasVec_6),
    .io_inConf_bits_confneuralNetsbiasVec_7(wellness_io_inConf_bits_confneuralNetsbiasVec_7),
    .io_inConf_bits_confneuralNetsbiasVec_8(wellness_io_inConf_bits_confneuralNetsbiasVec_8),
    .io_inConf_bits_confneuralNetsbiasVec_9(wellness_io_inConf_bits_confneuralNetsbiasVec_9),
    .io_inConf_bits_confneuralNetsbiasVec_10(wellness_io_inConf_bits_confneuralNetsbiasVec_10),
    .io_inConf_bits_confneuralNetsbiasVec_11(wellness_io_inConf_bits_confneuralNetsbiasVec_11),
    .io_inConf_bits_confneuralNetsbiasVec_12(wellness_io_inConf_bits_confneuralNetsbiasVec_12),
    .io_inConf_bits_confneuralNetsbiasVec_13(wellness_io_inConf_bits_confneuralNetsbiasVec_13),
    .io_inConf_bits_confneuralNetsbiasVec_14(wellness_io_inConf_bits_confneuralNetsbiasVec_14),
    .io_inConf_bits_confneuralNetsbiasVec_15(wellness_io_inConf_bits_confneuralNetsbiasVec_15),
    .io_inConf_bits_confneuralNetsbiasVec_16(wellness_io_inConf_bits_confneuralNetsbiasVec_16),
    .io_inConf_bits_confneuralNetsbiasVec_17(wellness_io_inConf_bits_confneuralNetsbiasVec_17),
    .io_inConf_bits_confneuralNetsbiasVec_18(wellness_io_inConf_bits_confneuralNetsbiasVec_18),
    .io_inConf_bits_confneuralNetsbiasVec_19(wellness_io_inConf_bits_confneuralNetsbiasVec_19),
    .io_inConf_bits_confneuralNetsbiasVec_20(wellness_io_inConf_bits_confneuralNetsbiasVec_20),
    .io_inConf_bits_confneuralNetsbiasVec_21(wellness_io_inConf_bits_confneuralNetsbiasVec_21),
    .io_inConf_bits_confneuralNetsbiasVec_22(wellness_io_inConf_bits_confneuralNetsbiasVec_22),
    .io_inConf_bits_confneuralNetsbiasVec_23(wellness_io_inConf_bits_confneuralNetsbiasVec_23),
    .io_inConf_bits_confneuralNetsbiasVec_24(wellness_io_inConf_bits_confneuralNetsbiasVec_24),
    .io_inConf_bits_confneuralNetsbiasVec_25(wellness_io_inConf_bits_confneuralNetsbiasVec_25),
    .io_inConf_bits_confneuralNetsbiasVec_26(wellness_io_inConf_bits_confneuralNetsbiasVec_26),
    .io_inConf_bits_confneuralNetsbiasVec_27(wellness_io_inConf_bits_confneuralNetsbiasVec_27),
    .io_inConf_bits_confneuralNetsbiasVec_28(wellness_io_inConf_bits_confneuralNetsbiasVec_28),
    .io_inConf_bits_confneuralNetsbiasVec_29(wellness_io_inConf_bits_confneuralNetsbiasVec_29),
    .io_inConf_bits_confneuralNetsbiasVec_30(wellness_io_inConf_bits_confneuralNetsbiasVec_30),
    .io_inConf_bits_confneuralNetsbiasVec_31(wellness_io_inConf_bits_confneuralNetsbiasVec_31),
    .io_inConf_bits_confneuralNetsbiasVec_32(wellness_io_inConf_bits_confneuralNetsbiasVec_32),
    .io_inConf_bits_confneuralNetsbiasVec_33(wellness_io_inConf_bits_confneuralNetsbiasVec_33),
    .io_inConf_bits_confneuralNetsbiasVec_34(wellness_io_inConf_bits_confneuralNetsbiasVec_34),
    .io_inConf_bits_confneuralNetsbiasVec_35(wellness_io_inConf_bits_confneuralNetsbiasVec_35),
    .io_inConf_bits_confneuralNetsbiasVec_36(wellness_io_inConf_bits_confneuralNetsbiasVec_36),
    .io_inConf_bits_confneuralNetsbiasVec_37(wellness_io_inConf_bits_confneuralNetsbiasVec_37),
    .io_inConf_bits_confneuralNetsbiasVec_38(wellness_io_inConf_bits_confneuralNetsbiasVec_38),
    .io_inConf_bits_confneuralNetsbiasVec_39(wellness_io_inConf_bits_confneuralNetsbiasVec_39),
    .io_inConf_bits_confneuralNetsbiasVec_40(wellness_io_inConf_bits_confneuralNetsbiasVec_40),
    .io_inConf_bits_confneuralNetsbiasVec_41(wellness_io_inConf_bits_confneuralNetsbiasVec_41),
    .io_inConf_bits_confneuralNetsbiasVec_42(wellness_io_inConf_bits_confneuralNetsbiasVec_42),
    .io_inConf_bits_confneuralNetsbiasVec_43(wellness_io_inConf_bits_confneuralNetsbiasVec_43),
    .io_inConf_bits_confneuralNetsbiasVec_44(wellness_io_inConf_bits_confneuralNetsbiasVec_44),
    .io_inConf_bits_confneuralNetsbiasVec_45(wellness_io_inConf_bits_confneuralNetsbiasVec_45),
    .io_inConf_bits_confneuralNetsbiasVec_46(wellness_io_inConf_bits_confneuralNetsbiasVec_46),
    .io_inConf_bits_confneuralNetsbiasVec_47(wellness_io_inConf_bits_confneuralNetsbiasVec_47),
    .io_inConf_bits_confneuralNetsbiasVec_48(wellness_io_inConf_bits_confneuralNetsbiasVec_48),
    .io_inConf_bits_confneuralNetsbiasVec_49(wellness_io_inConf_bits_confneuralNetsbiasVec_49),
    .io_inConf_bits_confneuralNetsbiasVec_50(wellness_io_inConf_bits_confneuralNetsbiasVec_50),
    .io_inConf_bits_confneuralNetsbiasVec_51(wellness_io_inConf_bits_confneuralNetsbiasVec_51),
    .io_inConf_bits_confneuralNetsbiasVec_52(wellness_io_inConf_bits_confneuralNetsbiasVec_52),
    .io_inConf_bits_confneuralNetsbiasVec_53(wellness_io_inConf_bits_confneuralNetsbiasVec_53),
    .io_inConf_bits_confneuralNetsbiasVec_54(wellness_io_inConf_bits_confneuralNetsbiasVec_54),
    .io_inConf_bits_confneuralNetsbiasVec_55(wellness_io_inConf_bits_confneuralNetsbiasVec_55),
    .io_inConf_bits_confneuralNetsbiasVec_56(wellness_io_inConf_bits_confneuralNetsbiasVec_56),
    .io_inConf_bits_confneuralNetsbiasVec_57(wellness_io_inConf_bits_confneuralNetsbiasVec_57),
    .io_inConf_bits_confneuralNetsbiasVec_58(wellness_io_inConf_bits_confneuralNetsbiasVec_58),
    .io_inConf_bits_confneuralNetsbiasVec_59(wellness_io_inConf_bits_confneuralNetsbiasVec_59),
    .io_inConf_bits_confneuralNetsbiasVec_60(wellness_io_inConf_bits_confneuralNetsbiasVec_60),
    .io_inConf_bits_confneuralNetsbiasVec_61(wellness_io_inConf_bits_confneuralNetsbiasVec_61),
    .io_inConf_bits_confneuralNetsbiasVec_62(wellness_io_inConf_bits_confneuralNetsbiasVec_62),
    .io_inConf_bits_confneuralNetsbiasVec_63(wellness_io_inConf_bits_confneuralNetsbiasVec_63),
    .io_inConf_bits_confneuralNetsbiasVec_64(wellness_io_inConf_bits_confneuralNetsbiasVec_64),
    .io_inConf_bits_confneuralNetsbiasVec_65(wellness_io_inConf_bits_confneuralNetsbiasVec_65),
    .io_inConf_bits_confneuralNetsbiasVec_66(wellness_io_inConf_bits_confneuralNetsbiasVec_66),
    .io_inConf_bits_confneuralNetsbiasVec_67(wellness_io_inConf_bits_confneuralNetsbiasVec_67),
    .io_inConf_bits_confneuralNetsbiasVec_68(wellness_io_inConf_bits_confneuralNetsbiasVec_68),
    .io_inConf_bits_confneuralNetsbiasVec_69(wellness_io_inConf_bits_confneuralNetsbiasVec_69),
    .io_inConf_bits_confneuralNetsbiasVec_70(wellness_io_inConf_bits_confneuralNetsbiasVec_70),
    .io_inConf_bits_confneuralNetsbiasVec_71(wellness_io_inConf_bits_confneuralNetsbiasVec_71),
    .io_inConf_bits_confneuralNetsbiasVec_72(wellness_io_inConf_bits_confneuralNetsbiasVec_72),
    .io_inConf_bits_confneuralNetsbiasVec_73(wellness_io_inConf_bits_confneuralNetsbiasVec_73),
    .io_inConf_bits_confneuralNetsbiasVec_74(wellness_io_inConf_bits_confneuralNetsbiasVec_74),
    .io_inConf_bits_confneuralNetsbiasVec_75(wellness_io_inConf_bits_confneuralNetsbiasVec_75),
    .io_inConf_bits_confneuralNetsbiasVec_76(wellness_io_inConf_bits_confneuralNetsbiasVec_76),
    .io_inConf_bits_confneuralNetsbiasVec_77(wellness_io_inConf_bits_confneuralNetsbiasVec_77),
    .io_inConf_bits_confneuralNetsbiasVec_78(wellness_io_inConf_bits_confneuralNetsbiasVec_78),
    .io_inConf_bits_confneuralNetsbiasVec_79(wellness_io_inConf_bits_confneuralNetsbiasVec_79),
    .io_inConf_bits_confneuralNetsbiasVec_80(wellness_io_inConf_bits_confneuralNetsbiasVec_80),
    .io_inConf_bits_confneuralNetsbiasVec_81(wellness_io_inConf_bits_confneuralNetsbiasVec_81),
    .io_inConf_bits_confneuralNetsbiasVec_82(wellness_io_inConf_bits_confneuralNetsbiasVec_82),
    .io_inConf_bits_confneuralNetsbiasVec_83(wellness_io_inConf_bits_confneuralNetsbiasVec_83),
    .io_inConf_bits_confneuralNetsbiasVec_84(wellness_io_inConf_bits_confneuralNetsbiasVec_84),
    .io_inConf_bits_confneuralNetsbiasVec_85(wellness_io_inConf_bits_confneuralNetsbiasVec_85),
    .io_inConf_bits_confneuralNetsbiasVec_86(wellness_io_inConf_bits_confneuralNetsbiasVec_86),
    .io_inConf_bits_confneuralNetsbiasVec_87(wellness_io_inConf_bits_confneuralNetsbiasVec_87),
    .io_inConf_bits_confneuralNetsbiasVec_88(wellness_io_inConf_bits_confneuralNetsbiasVec_88),
    .io_inConf_bits_confneuralNetsbiasVec_89(wellness_io_inConf_bits_confneuralNetsbiasVec_89),
    .io_inConf_bits_confneuralNetsbiasVec_90(wellness_io_inConf_bits_confneuralNetsbiasVec_90),
    .io_inConf_bits_confneuralNetsbiasVec_91(wellness_io_inConf_bits_confneuralNetsbiasVec_91),
    .io_inConf_bits_confneuralNetsbiasVec_92(wellness_io_inConf_bits_confneuralNetsbiasVec_92),
    .io_inConf_bits_confneuralNetsbiasVec_93(wellness_io_inConf_bits_confneuralNetsbiasVec_93),
    .io_inConf_bits_confneuralNetsbiasVec_94(wellness_io_inConf_bits_confneuralNetsbiasVec_94),
    .io_inConf_bits_confneuralNetsbiasVec_95(wellness_io_inConf_bits_confneuralNetsbiasVec_95),
    .io_inConf_bits_confneuralNetsbiasVec_96(wellness_io_inConf_bits_confneuralNetsbiasVec_96),
    .io_inConf_bits_confneuralNetsbiasVec_97(wellness_io_inConf_bits_confneuralNetsbiasVec_97),
    .io_inConf_bits_confneuralNetsbiasVec_98(wellness_io_inConf_bits_confneuralNetsbiasVec_98),
    .io_inConf_bits_confneuralNetsbiasVec_99(wellness_io_inConf_bits_confneuralNetsbiasVec_99),
    .io_inConf_bits_confneuralNetsbiasScalar_0(wellness_io_inConf_bits_confneuralNetsbiasScalar_0),
    .io_inConf_bits_confInputMuxSel(wellness_io_inConf_bits_confInputMuxSel),
    .io_out_valid(wellness_io_out_valid),
    .io_out_bits(wellness_io_out_bits),
    .io_rawVotes(wellness_io_rawVotes)
  );
  ConfigurationMemory configurationMemory ( // @[Wellness.scala 398:37]
    .clock(configurationMemory_clock),
    .reset(configurationMemory_reset),
    .io_in_valid(configurationMemory_io_in_valid),
    .io_in_bits_wrdata(configurationMemory_io_in_bits_wrdata),
    .io_in_bits_wraddr(configurationMemory_io_in_bits_wraddr),
    .io_out_bits_confneuralNetsweightMatrix_0_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_0_0),
    .io_out_bits_confneuralNetsweightMatrix_0_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_0_1),
    .io_out_bits_confneuralNetsweightMatrix_0_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_0_2),
    .io_out_bits_confneuralNetsweightMatrix_0_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_0_3),
    .io_out_bits_confneuralNetsweightMatrix_1_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_1_0),
    .io_out_bits_confneuralNetsweightMatrix_1_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_1_1),
    .io_out_bits_confneuralNetsweightMatrix_1_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_1_2),
    .io_out_bits_confneuralNetsweightMatrix_1_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_1_3),
    .io_out_bits_confneuralNetsweightMatrix_2_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_2_0),
    .io_out_bits_confneuralNetsweightMatrix_2_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_2_1),
    .io_out_bits_confneuralNetsweightMatrix_2_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_2_2),
    .io_out_bits_confneuralNetsweightMatrix_2_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_2_3),
    .io_out_bits_confneuralNetsweightMatrix_3_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_3_0),
    .io_out_bits_confneuralNetsweightMatrix_3_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_3_1),
    .io_out_bits_confneuralNetsweightMatrix_3_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_3_2),
    .io_out_bits_confneuralNetsweightMatrix_3_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_3_3),
    .io_out_bits_confneuralNetsweightMatrix_4_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_4_0),
    .io_out_bits_confneuralNetsweightMatrix_4_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_4_1),
    .io_out_bits_confneuralNetsweightMatrix_4_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_4_2),
    .io_out_bits_confneuralNetsweightMatrix_4_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_4_3),
    .io_out_bits_confneuralNetsweightMatrix_5_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_5_0),
    .io_out_bits_confneuralNetsweightMatrix_5_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_5_1),
    .io_out_bits_confneuralNetsweightMatrix_5_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_5_2),
    .io_out_bits_confneuralNetsweightMatrix_5_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_5_3),
    .io_out_bits_confneuralNetsweightMatrix_6_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_6_0),
    .io_out_bits_confneuralNetsweightMatrix_6_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_6_1),
    .io_out_bits_confneuralNetsweightMatrix_6_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_6_2),
    .io_out_bits_confneuralNetsweightMatrix_6_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_6_3),
    .io_out_bits_confneuralNetsweightMatrix_7_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_7_0),
    .io_out_bits_confneuralNetsweightMatrix_7_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_7_1),
    .io_out_bits_confneuralNetsweightMatrix_7_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_7_2),
    .io_out_bits_confneuralNetsweightMatrix_7_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_7_3),
    .io_out_bits_confneuralNetsweightMatrix_8_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_8_0),
    .io_out_bits_confneuralNetsweightMatrix_8_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_8_1),
    .io_out_bits_confneuralNetsweightMatrix_8_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_8_2),
    .io_out_bits_confneuralNetsweightMatrix_8_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_8_3),
    .io_out_bits_confneuralNetsweightMatrix_9_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_9_0),
    .io_out_bits_confneuralNetsweightMatrix_9_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_9_1),
    .io_out_bits_confneuralNetsweightMatrix_9_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_9_2),
    .io_out_bits_confneuralNetsweightMatrix_9_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_9_3),
    .io_out_bits_confneuralNetsweightMatrix_10_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_10_0),
    .io_out_bits_confneuralNetsweightMatrix_10_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_10_1),
    .io_out_bits_confneuralNetsweightMatrix_10_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_10_2),
    .io_out_bits_confneuralNetsweightMatrix_10_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_10_3),
    .io_out_bits_confneuralNetsweightMatrix_11_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_11_0),
    .io_out_bits_confneuralNetsweightMatrix_11_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_11_1),
    .io_out_bits_confneuralNetsweightMatrix_11_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_11_2),
    .io_out_bits_confneuralNetsweightMatrix_11_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_11_3),
    .io_out_bits_confneuralNetsweightMatrix_12_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_12_0),
    .io_out_bits_confneuralNetsweightMatrix_12_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_12_1),
    .io_out_bits_confneuralNetsweightMatrix_12_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_12_2),
    .io_out_bits_confneuralNetsweightMatrix_12_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_12_3),
    .io_out_bits_confneuralNetsweightMatrix_13_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_13_0),
    .io_out_bits_confneuralNetsweightMatrix_13_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_13_1),
    .io_out_bits_confneuralNetsweightMatrix_13_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_13_2),
    .io_out_bits_confneuralNetsweightMatrix_13_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_13_3),
    .io_out_bits_confneuralNetsweightMatrix_14_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_14_0),
    .io_out_bits_confneuralNetsweightMatrix_14_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_14_1),
    .io_out_bits_confneuralNetsweightMatrix_14_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_14_2),
    .io_out_bits_confneuralNetsweightMatrix_14_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_14_3),
    .io_out_bits_confneuralNetsweightMatrix_15_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_15_0),
    .io_out_bits_confneuralNetsweightMatrix_15_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_15_1),
    .io_out_bits_confneuralNetsweightMatrix_15_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_15_2),
    .io_out_bits_confneuralNetsweightMatrix_15_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_15_3),
    .io_out_bits_confneuralNetsweightMatrix_16_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_16_0),
    .io_out_bits_confneuralNetsweightMatrix_16_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_16_1),
    .io_out_bits_confneuralNetsweightMatrix_16_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_16_2),
    .io_out_bits_confneuralNetsweightMatrix_16_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_16_3),
    .io_out_bits_confneuralNetsweightMatrix_17_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_17_0),
    .io_out_bits_confneuralNetsweightMatrix_17_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_17_1),
    .io_out_bits_confneuralNetsweightMatrix_17_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_17_2),
    .io_out_bits_confneuralNetsweightMatrix_17_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_17_3),
    .io_out_bits_confneuralNetsweightMatrix_18_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_18_0),
    .io_out_bits_confneuralNetsweightMatrix_18_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_18_1),
    .io_out_bits_confneuralNetsweightMatrix_18_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_18_2),
    .io_out_bits_confneuralNetsweightMatrix_18_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_18_3),
    .io_out_bits_confneuralNetsweightMatrix_19_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_19_0),
    .io_out_bits_confneuralNetsweightMatrix_19_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_19_1),
    .io_out_bits_confneuralNetsweightMatrix_19_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_19_2),
    .io_out_bits_confneuralNetsweightMatrix_19_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_19_3),
    .io_out_bits_confneuralNetsweightMatrix_20_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_20_0),
    .io_out_bits_confneuralNetsweightMatrix_20_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_20_1),
    .io_out_bits_confneuralNetsweightMatrix_20_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_20_2),
    .io_out_bits_confneuralNetsweightMatrix_20_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_20_3),
    .io_out_bits_confneuralNetsweightMatrix_21_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_21_0),
    .io_out_bits_confneuralNetsweightMatrix_21_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_21_1),
    .io_out_bits_confneuralNetsweightMatrix_21_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_21_2),
    .io_out_bits_confneuralNetsweightMatrix_21_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_21_3),
    .io_out_bits_confneuralNetsweightMatrix_22_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_22_0),
    .io_out_bits_confneuralNetsweightMatrix_22_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_22_1),
    .io_out_bits_confneuralNetsweightMatrix_22_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_22_2),
    .io_out_bits_confneuralNetsweightMatrix_22_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_22_3),
    .io_out_bits_confneuralNetsweightMatrix_23_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_23_0),
    .io_out_bits_confneuralNetsweightMatrix_23_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_23_1),
    .io_out_bits_confneuralNetsweightMatrix_23_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_23_2),
    .io_out_bits_confneuralNetsweightMatrix_23_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_23_3),
    .io_out_bits_confneuralNetsweightMatrix_24_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_24_0),
    .io_out_bits_confneuralNetsweightMatrix_24_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_24_1),
    .io_out_bits_confneuralNetsweightMatrix_24_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_24_2),
    .io_out_bits_confneuralNetsweightMatrix_24_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_24_3),
    .io_out_bits_confneuralNetsweightMatrix_25_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_25_0),
    .io_out_bits_confneuralNetsweightMatrix_25_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_25_1),
    .io_out_bits_confneuralNetsweightMatrix_25_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_25_2),
    .io_out_bits_confneuralNetsweightMatrix_25_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_25_3),
    .io_out_bits_confneuralNetsweightMatrix_26_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_26_0),
    .io_out_bits_confneuralNetsweightMatrix_26_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_26_1),
    .io_out_bits_confneuralNetsweightMatrix_26_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_26_2),
    .io_out_bits_confneuralNetsweightMatrix_26_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_26_3),
    .io_out_bits_confneuralNetsweightMatrix_27_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_27_0),
    .io_out_bits_confneuralNetsweightMatrix_27_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_27_1),
    .io_out_bits_confneuralNetsweightMatrix_27_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_27_2),
    .io_out_bits_confneuralNetsweightMatrix_27_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_27_3),
    .io_out_bits_confneuralNetsweightMatrix_28_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_28_0),
    .io_out_bits_confneuralNetsweightMatrix_28_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_28_1),
    .io_out_bits_confneuralNetsweightMatrix_28_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_28_2),
    .io_out_bits_confneuralNetsweightMatrix_28_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_28_3),
    .io_out_bits_confneuralNetsweightMatrix_29_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_29_0),
    .io_out_bits_confneuralNetsweightMatrix_29_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_29_1),
    .io_out_bits_confneuralNetsweightMatrix_29_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_29_2),
    .io_out_bits_confneuralNetsweightMatrix_29_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_29_3),
    .io_out_bits_confneuralNetsweightMatrix_30_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_30_0),
    .io_out_bits_confneuralNetsweightMatrix_30_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_30_1),
    .io_out_bits_confneuralNetsweightMatrix_30_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_30_2),
    .io_out_bits_confneuralNetsweightMatrix_30_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_30_3),
    .io_out_bits_confneuralNetsweightMatrix_31_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_31_0),
    .io_out_bits_confneuralNetsweightMatrix_31_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_31_1),
    .io_out_bits_confneuralNetsweightMatrix_31_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_31_2),
    .io_out_bits_confneuralNetsweightMatrix_31_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_31_3),
    .io_out_bits_confneuralNetsweightMatrix_32_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_32_0),
    .io_out_bits_confneuralNetsweightMatrix_32_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_32_1),
    .io_out_bits_confneuralNetsweightMatrix_32_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_32_2),
    .io_out_bits_confneuralNetsweightMatrix_32_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_32_3),
    .io_out_bits_confneuralNetsweightMatrix_33_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_33_0),
    .io_out_bits_confneuralNetsweightMatrix_33_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_33_1),
    .io_out_bits_confneuralNetsweightMatrix_33_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_33_2),
    .io_out_bits_confneuralNetsweightMatrix_33_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_33_3),
    .io_out_bits_confneuralNetsweightMatrix_34_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_34_0),
    .io_out_bits_confneuralNetsweightMatrix_34_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_34_1),
    .io_out_bits_confneuralNetsweightMatrix_34_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_34_2),
    .io_out_bits_confneuralNetsweightMatrix_34_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_34_3),
    .io_out_bits_confneuralNetsweightMatrix_35_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_35_0),
    .io_out_bits_confneuralNetsweightMatrix_35_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_35_1),
    .io_out_bits_confneuralNetsweightMatrix_35_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_35_2),
    .io_out_bits_confneuralNetsweightMatrix_35_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_35_3),
    .io_out_bits_confneuralNetsweightMatrix_36_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_36_0),
    .io_out_bits_confneuralNetsweightMatrix_36_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_36_1),
    .io_out_bits_confneuralNetsweightMatrix_36_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_36_2),
    .io_out_bits_confneuralNetsweightMatrix_36_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_36_3),
    .io_out_bits_confneuralNetsweightMatrix_37_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_37_0),
    .io_out_bits_confneuralNetsweightMatrix_37_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_37_1),
    .io_out_bits_confneuralNetsweightMatrix_37_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_37_2),
    .io_out_bits_confneuralNetsweightMatrix_37_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_37_3),
    .io_out_bits_confneuralNetsweightMatrix_38_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_38_0),
    .io_out_bits_confneuralNetsweightMatrix_38_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_38_1),
    .io_out_bits_confneuralNetsweightMatrix_38_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_38_2),
    .io_out_bits_confneuralNetsweightMatrix_38_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_38_3),
    .io_out_bits_confneuralNetsweightMatrix_39_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_39_0),
    .io_out_bits_confneuralNetsweightMatrix_39_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_39_1),
    .io_out_bits_confneuralNetsweightMatrix_39_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_39_2),
    .io_out_bits_confneuralNetsweightMatrix_39_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_39_3),
    .io_out_bits_confneuralNetsweightMatrix_40_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_40_0),
    .io_out_bits_confneuralNetsweightMatrix_40_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_40_1),
    .io_out_bits_confneuralNetsweightMatrix_40_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_40_2),
    .io_out_bits_confneuralNetsweightMatrix_40_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_40_3),
    .io_out_bits_confneuralNetsweightMatrix_41_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_41_0),
    .io_out_bits_confneuralNetsweightMatrix_41_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_41_1),
    .io_out_bits_confneuralNetsweightMatrix_41_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_41_2),
    .io_out_bits_confneuralNetsweightMatrix_41_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_41_3),
    .io_out_bits_confneuralNetsweightMatrix_42_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_42_0),
    .io_out_bits_confneuralNetsweightMatrix_42_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_42_1),
    .io_out_bits_confneuralNetsweightMatrix_42_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_42_2),
    .io_out_bits_confneuralNetsweightMatrix_42_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_42_3),
    .io_out_bits_confneuralNetsweightMatrix_43_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_43_0),
    .io_out_bits_confneuralNetsweightMatrix_43_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_43_1),
    .io_out_bits_confneuralNetsweightMatrix_43_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_43_2),
    .io_out_bits_confneuralNetsweightMatrix_43_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_43_3),
    .io_out_bits_confneuralNetsweightMatrix_44_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_44_0),
    .io_out_bits_confneuralNetsweightMatrix_44_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_44_1),
    .io_out_bits_confneuralNetsweightMatrix_44_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_44_2),
    .io_out_bits_confneuralNetsweightMatrix_44_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_44_3),
    .io_out_bits_confneuralNetsweightMatrix_45_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_45_0),
    .io_out_bits_confneuralNetsweightMatrix_45_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_45_1),
    .io_out_bits_confneuralNetsweightMatrix_45_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_45_2),
    .io_out_bits_confneuralNetsweightMatrix_45_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_45_3),
    .io_out_bits_confneuralNetsweightMatrix_46_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_46_0),
    .io_out_bits_confneuralNetsweightMatrix_46_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_46_1),
    .io_out_bits_confneuralNetsweightMatrix_46_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_46_2),
    .io_out_bits_confneuralNetsweightMatrix_46_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_46_3),
    .io_out_bits_confneuralNetsweightMatrix_47_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_47_0),
    .io_out_bits_confneuralNetsweightMatrix_47_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_47_1),
    .io_out_bits_confneuralNetsweightMatrix_47_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_47_2),
    .io_out_bits_confneuralNetsweightMatrix_47_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_47_3),
    .io_out_bits_confneuralNetsweightMatrix_48_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_48_0),
    .io_out_bits_confneuralNetsweightMatrix_48_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_48_1),
    .io_out_bits_confneuralNetsweightMatrix_48_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_48_2),
    .io_out_bits_confneuralNetsweightMatrix_48_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_48_3),
    .io_out_bits_confneuralNetsweightMatrix_49_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_49_0),
    .io_out_bits_confneuralNetsweightMatrix_49_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_49_1),
    .io_out_bits_confneuralNetsweightMatrix_49_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_49_2),
    .io_out_bits_confneuralNetsweightMatrix_49_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_49_3),
    .io_out_bits_confneuralNetsweightMatrix_50_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_50_0),
    .io_out_bits_confneuralNetsweightMatrix_50_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_50_1),
    .io_out_bits_confneuralNetsweightMatrix_50_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_50_2),
    .io_out_bits_confneuralNetsweightMatrix_50_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_50_3),
    .io_out_bits_confneuralNetsweightMatrix_51_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_51_0),
    .io_out_bits_confneuralNetsweightMatrix_51_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_51_1),
    .io_out_bits_confneuralNetsweightMatrix_51_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_51_2),
    .io_out_bits_confneuralNetsweightMatrix_51_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_51_3),
    .io_out_bits_confneuralNetsweightMatrix_52_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_52_0),
    .io_out_bits_confneuralNetsweightMatrix_52_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_52_1),
    .io_out_bits_confneuralNetsweightMatrix_52_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_52_2),
    .io_out_bits_confneuralNetsweightMatrix_52_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_52_3),
    .io_out_bits_confneuralNetsweightMatrix_53_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_53_0),
    .io_out_bits_confneuralNetsweightMatrix_53_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_53_1),
    .io_out_bits_confneuralNetsweightMatrix_53_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_53_2),
    .io_out_bits_confneuralNetsweightMatrix_53_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_53_3),
    .io_out_bits_confneuralNetsweightMatrix_54_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_54_0),
    .io_out_bits_confneuralNetsweightMatrix_54_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_54_1),
    .io_out_bits_confneuralNetsweightMatrix_54_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_54_2),
    .io_out_bits_confneuralNetsweightMatrix_54_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_54_3),
    .io_out_bits_confneuralNetsweightMatrix_55_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_55_0),
    .io_out_bits_confneuralNetsweightMatrix_55_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_55_1),
    .io_out_bits_confneuralNetsweightMatrix_55_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_55_2),
    .io_out_bits_confneuralNetsweightMatrix_55_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_55_3),
    .io_out_bits_confneuralNetsweightMatrix_56_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_56_0),
    .io_out_bits_confneuralNetsweightMatrix_56_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_56_1),
    .io_out_bits_confneuralNetsweightMatrix_56_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_56_2),
    .io_out_bits_confneuralNetsweightMatrix_56_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_56_3),
    .io_out_bits_confneuralNetsweightMatrix_57_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_57_0),
    .io_out_bits_confneuralNetsweightMatrix_57_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_57_1),
    .io_out_bits_confneuralNetsweightMatrix_57_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_57_2),
    .io_out_bits_confneuralNetsweightMatrix_57_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_57_3),
    .io_out_bits_confneuralNetsweightMatrix_58_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_58_0),
    .io_out_bits_confneuralNetsweightMatrix_58_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_58_1),
    .io_out_bits_confneuralNetsweightMatrix_58_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_58_2),
    .io_out_bits_confneuralNetsweightMatrix_58_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_58_3),
    .io_out_bits_confneuralNetsweightMatrix_59_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_59_0),
    .io_out_bits_confneuralNetsweightMatrix_59_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_59_1),
    .io_out_bits_confneuralNetsweightMatrix_59_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_59_2),
    .io_out_bits_confneuralNetsweightMatrix_59_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_59_3),
    .io_out_bits_confneuralNetsweightMatrix_60_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_60_0),
    .io_out_bits_confneuralNetsweightMatrix_60_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_60_1),
    .io_out_bits_confneuralNetsweightMatrix_60_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_60_2),
    .io_out_bits_confneuralNetsweightMatrix_60_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_60_3),
    .io_out_bits_confneuralNetsweightMatrix_61_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_61_0),
    .io_out_bits_confneuralNetsweightMatrix_61_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_61_1),
    .io_out_bits_confneuralNetsweightMatrix_61_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_61_2),
    .io_out_bits_confneuralNetsweightMatrix_61_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_61_3),
    .io_out_bits_confneuralNetsweightMatrix_62_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_62_0),
    .io_out_bits_confneuralNetsweightMatrix_62_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_62_1),
    .io_out_bits_confneuralNetsweightMatrix_62_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_62_2),
    .io_out_bits_confneuralNetsweightMatrix_62_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_62_3),
    .io_out_bits_confneuralNetsweightMatrix_63_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_63_0),
    .io_out_bits_confneuralNetsweightMatrix_63_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_63_1),
    .io_out_bits_confneuralNetsweightMatrix_63_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_63_2),
    .io_out_bits_confneuralNetsweightMatrix_63_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_63_3),
    .io_out_bits_confneuralNetsweightMatrix_64_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_64_0),
    .io_out_bits_confneuralNetsweightMatrix_64_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_64_1),
    .io_out_bits_confneuralNetsweightMatrix_64_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_64_2),
    .io_out_bits_confneuralNetsweightMatrix_64_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_64_3),
    .io_out_bits_confneuralNetsweightMatrix_65_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_65_0),
    .io_out_bits_confneuralNetsweightMatrix_65_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_65_1),
    .io_out_bits_confneuralNetsweightMatrix_65_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_65_2),
    .io_out_bits_confneuralNetsweightMatrix_65_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_65_3),
    .io_out_bits_confneuralNetsweightMatrix_66_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_66_0),
    .io_out_bits_confneuralNetsweightMatrix_66_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_66_1),
    .io_out_bits_confneuralNetsweightMatrix_66_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_66_2),
    .io_out_bits_confneuralNetsweightMatrix_66_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_66_3),
    .io_out_bits_confneuralNetsweightMatrix_67_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_67_0),
    .io_out_bits_confneuralNetsweightMatrix_67_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_67_1),
    .io_out_bits_confneuralNetsweightMatrix_67_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_67_2),
    .io_out_bits_confneuralNetsweightMatrix_67_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_67_3),
    .io_out_bits_confneuralNetsweightMatrix_68_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_68_0),
    .io_out_bits_confneuralNetsweightMatrix_68_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_68_1),
    .io_out_bits_confneuralNetsweightMatrix_68_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_68_2),
    .io_out_bits_confneuralNetsweightMatrix_68_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_68_3),
    .io_out_bits_confneuralNetsweightMatrix_69_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_69_0),
    .io_out_bits_confneuralNetsweightMatrix_69_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_69_1),
    .io_out_bits_confneuralNetsweightMatrix_69_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_69_2),
    .io_out_bits_confneuralNetsweightMatrix_69_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_69_3),
    .io_out_bits_confneuralNetsweightMatrix_70_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_70_0),
    .io_out_bits_confneuralNetsweightMatrix_70_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_70_1),
    .io_out_bits_confneuralNetsweightMatrix_70_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_70_2),
    .io_out_bits_confneuralNetsweightMatrix_70_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_70_3),
    .io_out_bits_confneuralNetsweightMatrix_71_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_71_0),
    .io_out_bits_confneuralNetsweightMatrix_71_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_71_1),
    .io_out_bits_confneuralNetsweightMatrix_71_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_71_2),
    .io_out_bits_confneuralNetsweightMatrix_71_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_71_3),
    .io_out_bits_confneuralNetsweightMatrix_72_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_72_0),
    .io_out_bits_confneuralNetsweightMatrix_72_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_72_1),
    .io_out_bits_confneuralNetsweightMatrix_72_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_72_2),
    .io_out_bits_confneuralNetsweightMatrix_72_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_72_3),
    .io_out_bits_confneuralNetsweightMatrix_73_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_73_0),
    .io_out_bits_confneuralNetsweightMatrix_73_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_73_1),
    .io_out_bits_confneuralNetsweightMatrix_73_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_73_2),
    .io_out_bits_confneuralNetsweightMatrix_73_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_73_3),
    .io_out_bits_confneuralNetsweightMatrix_74_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_74_0),
    .io_out_bits_confneuralNetsweightMatrix_74_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_74_1),
    .io_out_bits_confneuralNetsweightMatrix_74_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_74_2),
    .io_out_bits_confneuralNetsweightMatrix_74_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_74_3),
    .io_out_bits_confneuralNetsweightMatrix_75_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_75_0),
    .io_out_bits_confneuralNetsweightMatrix_75_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_75_1),
    .io_out_bits_confneuralNetsweightMatrix_75_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_75_2),
    .io_out_bits_confneuralNetsweightMatrix_75_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_75_3),
    .io_out_bits_confneuralNetsweightMatrix_76_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_76_0),
    .io_out_bits_confneuralNetsweightMatrix_76_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_76_1),
    .io_out_bits_confneuralNetsweightMatrix_76_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_76_2),
    .io_out_bits_confneuralNetsweightMatrix_76_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_76_3),
    .io_out_bits_confneuralNetsweightMatrix_77_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_77_0),
    .io_out_bits_confneuralNetsweightMatrix_77_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_77_1),
    .io_out_bits_confneuralNetsweightMatrix_77_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_77_2),
    .io_out_bits_confneuralNetsweightMatrix_77_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_77_3),
    .io_out_bits_confneuralNetsweightMatrix_78_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_78_0),
    .io_out_bits_confneuralNetsweightMatrix_78_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_78_1),
    .io_out_bits_confneuralNetsweightMatrix_78_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_78_2),
    .io_out_bits_confneuralNetsweightMatrix_78_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_78_3),
    .io_out_bits_confneuralNetsweightMatrix_79_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_79_0),
    .io_out_bits_confneuralNetsweightMatrix_79_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_79_1),
    .io_out_bits_confneuralNetsweightMatrix_79_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_79_2),
    .io_out_bits_confneuralNetsweightMatrix_79_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_79_3),
    .io_out_bits_confneuralNetsweightMatrix_80_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_80_0),
    .io_out_bits_confneuralNetsweightMatrix_80_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_80_1),
    .io_out_bits_confneuralNetsweightMatrix_80_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_80_2),
    .io_out_bits_confneuralNetsweightMatrix_80_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_80_3),
    .io_out_bits_confneuralNetsweightMatrix_81_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_81_0),
    .io_out_bits_confneuralNetsweightMatrix_81_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_81_1),
    .io_out_bits_confneuralNetsweightMatrix_81_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_81_2),
    .io_out_bits_confneuralNetsweightMatrix_81_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_81_3),
    .io_out_bits_confneuralNetsweightMatrix_82_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_82_0),
    .io_out_bits_confneuralNetsweightMatrix_82_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_82_1),
    .io_out_bits_confneuralNetsweightMatrix_82_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_82_2),
    .io_out_bits_confneuralNetsweightMatrix_82_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_82_3),
    .io_out_bits_confneuralNetsweightMatrix_83_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_83_0),
    .io_out_bits_confneuralNetsweightMatrix_83_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_83_1),
    .io_out_bits_confneuralNetsweightMatrix_83_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_83_2),
    .io_out_bits_confneuralNetsweightMatrix_83_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_83_3),
    .io_out_bits_confneuralNetsweightMatrix_84_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_84_0),
    .io_out_bits_confneuralNetsweightMatrix_84_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_84_1),
    .io_out_bits_confneuralNetsweightMatrix_84_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_84_2),
    .io_out_bits_confneuralNetsweightMatrix_84_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_84_3),
    .io_out_bits_confneuralNetsweightMatrix_85_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_85_0),
    .io_out_bits_confneuralNetsweightMatrix_85_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_85_1),
    .io_out_bits_confneuralNetsweightMatrix_85_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_85_2),
    .io_out_bits_confneuralNetsweightMatrix_85_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_85_3),
    .io_out_bits_confneuralNetsweightMatrix_86_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_86_0),
    .io_out_bits_confneuralNetsweightMatrix_86_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_86_1),
    .io_out_bits_confneuralNetsweightMatrix_86_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_86_2),
    .io_out_bits_confneuralNetsweightMatrix_86_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_86_3),
    .io_out_bits_confneuralNetsweightMatrix_87_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_87_0),
    .io_out_bits_confneuralNetsweightMatrix_87_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_87_1),
    .io_out_bits_confneuralNetsweightMatrix_87_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_87_2),
    .io_out_bits_confneuralNetsweightMatrix_87_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_87_3),
    .io_out_bits_confneuralNetsweightMatrix_88_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_88_0),
    .io_out_bits_confneuralNetsweightMatrix_88_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_88_1),
    .io_out_bits_confneuralNetsweightMatrix_88_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_88_2),
    .io_out_bits_confneuralNetsweightMatrix_88_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_88_3),
    .io_out_bits_confneuralNetsweightMatrix_89_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_89_0),
    .io_out_bits_confneuralNetsweightMatrix_89_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_89_1),
    .io_out_bits_confneuralNetsweightMatrix_89_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_89_2),
    .io_out_bits_confneuralNetsweightMatrix_89_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_89_3),
    .io_out_bits_confneuralNetsweightMatrix_90_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_90_0),
    .io_out_bits_confneuralNetsweightMatrix_90_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_90_1),
    .io_out_bits_confneuralNetsweightMatrix_90_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_90_2),
    .io_out_bits_confneuralNetsweightMatrix_90_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_90_3),
    .io_out_bits_confneuralNetsweightMatrix_91_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_91_0),
    .io_out_bits_confneuralNetsweightMatrix_91_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_91_1),
    .io_out_bits_confneuralNetsweightMatrix_91_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_91_2),
    .io_out_bits_confneuralNetsweightMatrix_91_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_91_3),
    .io_out_bits_confneuralNetsweightMatrix_92_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_92_0),
    .io_out_bits_confneuralNetsweightMatrix_92_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_92_1),
    .io_out_bits_confneuralNetsweightMatrix_92_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_92_2),
    .io_out_bits_confneuralNetsweightMatrix_92_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_92_3),
    .io_out_bits_confneuralNetsweightMatrix_93_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_93_0),
    .io_out_bits_confneuralNetsweightMatrix_93_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_93_1),
    .io_out_bits_confneuralNetsweightMatrix_93_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_93_2),
    .io_out_bits_confneuralNetsweightMatrix_93_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_93_3),
    .io_out_bits_confneuralNetsweightMatrix_94_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_94_0),
    .io_out_bits_confneuralNetsweightMatrix_94_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_94_1),
    .io_out_bits_confneuralNetsweightMatrix_94_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_94_2),
    .io_out_bits_confneuralNetsweightMatrix_94_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_94_3),
    .io_out_bits_confneuralNetsweightMatrix_95_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_95_0),
    .io_out_bits_confneuralNetsweightMatrix_95_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_95_1),
    .io_out_bits_confneuralNetsweightMatrix_95_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_95_2),
    .io_out_bits_confneuralNetsweightMatrix_95_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_95_3),
    .io_out_bits_confneuralNetsweightMatrix_96_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_96_0),
    .io_out_bits_confneuralNetsweightMatrix_96_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_96_1),
    .io_out_bits_confneuralNetsweightMatrix_96_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_96_2),
    .io_out_bits_confneuralNetsweightMatrix_96_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_96_3),
    .io_out_bits_confneuralNetsweightMatrix_97_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_97_0),
    .io_out_bits_confneuralNetsweightMatrix_97_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_97_1),
    .io_out_bits_confneuralNetsweightMatrix_97_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_97_2),
    .io_out_bits_confneuralNetsweightMatrix_97_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_97_3),
    .io_out_bits_confneuralNetsweightMatrix_98_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_98_0),
    .io_out_bits_confneuralNetsweightMatrix_98_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_98_1),
    .io_out_bits_confneuralNetsweightMatrix_98_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_98_2),
    .io_out_bits_confneuralNetsweightMatrix_98_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_98_3),
    .io_out_bits_confneuralNetsweightMatrix_99_0(configurationMemory_io_out_bits_confneuralNetsweightMatrix_99_0),
    .io_out_bits_confneuralNetsweightMatrix_99_1(configurationMemory_io_out_bits_confneuralNetsweightMatrix_99_1),
    .io_out_bits_confneuralNetsweightMatrix_99_2(configurationMemory_io_out_bits_confneuralNetsweightMatrix_99_2),
    .io_out_bits_confneuralNetsweightMatrix_99_3(configurationMemory_io_out_bits_confneuralNetsweightMatrix_99_3),
    .io_out_bits_confneuralNetsweightVec_0(configurationMemory_io_out_bits_confneuralNetsweightVec_0),
    .io_out_bits_confneuralNetsweightVec_1(configurationMemory_io_out_bits_confneuralNetsweightVec_1),
    .io_out_bits_confneuralNetsweightVec_2(configurationMemory_io_out_bits_confneuralNetsweightVec_2),
    .io_out_bits_confneuralNetsweightVec_3(configurationMemory_io_out_bits_confneuralNetsweightVec_3),
    .io_out_bits_confneuralNetsweightVec_4(configurationMemory_io_out_bits_confneuralNetsweightVec_4),
    .io_out_bits_confneuralNetsweightVec_5(configurationMemory_io_out_bits_confneuralNetsweightVec_5),
    .io_out_bits_confneuralNetsweightVec_6(configurationMemory_io_out_bits_confneuralNetsweightVec_6),
    .io_out_bits_confneuralNetsweightVec_7(configurationMemory_io_out_bits_confneuralNetsweightVec_7),
    .io_out_bits_confneuralNetsweightVec_8(configurationMemory_io_out_bits_confneuralNetsweightVec_8),
    .io_out_bits_confneuralNetsweightVec_9(configurationMemory_io_out_bits_confneuralNetsweightVec_9),
    .io_out_bits_confneuralNetsweightVec_10(configurationMemory_io_out_bits_confneuralNetsweightVec_10),
    .io_out_bits_confneuralNetsweightVec_11(configurationMemory_io_out_bits_confneuralNetsweightVec_11),
    .io_out_bits_confneuralNetsweightVec_12(configurationMemory_io_out_bits_confneuralNetsweightVec_12),
    .io_out_bits_confneuralNetsweightVec_13(configurationMemory_io_out_bits_confneuralNetsweightVec_13),
    .io_out_bits_confneuralNetsweightVec_14(configurationMemory_io_out_bits_confneuralNetsweightVec_14),
    .io_out_bits_confneuralNetsweightVec_15(configurationMemory_io_out_bits_confneuralNetsweightVec_15),
    .io_out_bits_confneuralNetsweightVec_16(configurationMemory_io_out_bits_confneuralNetsweightVec_16),
    .io_out_bits_confneuralNetsweightVec_17(configurationMemory_io_out_bits_confneuralNetsweightVec_17),
    .io_out_bits_confneuralNetsweightVec_18(configurationMemory_io_out_bits_confneuralNetsweightVec_18),
    .io_out_bits_confneuralNetsweightVec_19(configurationMemory_io_out_bits_confneuralNetsweightVec_19),
    .io_out_bits_confneuralNetsweightVec_20(configurationMemory_io_out_bits_confneuralNetsweightVec_20),
    .io_out_bits_confneuralNetsweightVec_21(configurationMemory_io_out_bits_confneuralNetsweightVec_21),
    .io_out_bits_confneuralNetsweightVec_22(configurationMemory_io_out_bits_confneuralNetsweightVec_22),
    .io_out_bits_confneuralNetsweightVec_23(configurationMemory_io_out_bits_confneuralNetsweightVec_23),
    .io_out_bits_confneuralNetsweightVec_24(configurationMemory_io_out_bits_confneuralNetsweightVec_24),
    .io_out_bits_confneuralNetsweightVec_25(configurationMemory_io_out_bits_confneuralNetsweightVec_25),
    .io_out_bits_confneuralNetsweightVec_26(configurationMemory_io_out_bits_confneuralNetsweightVec_26),
    .io_out_bits_confneuralNetsweightVec_27(configurationMemory_io_out_bits_confneuralNetsweightVec_27),
    .io_out_bits_confneuralNetsweightVec_28(configurationMemory_io_out_bits_confneuralNetsweightVec_28),
    .io_out_bits_confneuralNetsweightVec_29(configurationMemory_io_out_bits_confneuralNetsweightVec_29),
    .io_out_bits_confneuralNetsweightVec_30(configurationMemory_io_out_bits_confneuralNetsweightVec_30),
    .io_out_bits_confneuralNetsweightVec_31(configurationMemory_io_out_bits_confneuralNetsweightVec_31),
    .io_out_bits_confneuralNetsweightVec_32(configurationMemory_io_out_bits_confneuralNetsweightVec_32),
    .io_out_bits_confneuralNetsweightVec_33(configurationMemory_io_out_bits_confneuralNetsweightVec_33),
    .io_out_bits_confneuralNetsweightVec_34(configurationMemory_io_out_bits_confneuralNetsweightVec_34),
    .io_out_bits_confneuralNetsweightVec_35(configurationMemory_io_out_bits_confneuralNetsweightVec_35),
    .io_out_bits_confneuralNetsweightVec_36(configurationMemory_io_out_bits_confneuralNetsweightVec_36),
    .io_out_bits_confneuralNetsweightVec_37(configurationMemory_io_out_bits_confneuralNetsweightVec_37),
    .io_out_bits_confneuralNetsweightVec_38(configurationMemory_io_out_bits_confneuralNetsweightVec_38),
    .io_out_bits_confneuralNetsweightVec_39(configurationMemory_io_out_bits_confneuralNetsweightVec_39),
    .io_out_bits_confneuralNetsweightVec_40(configurationMemory_io_out_bits_confneuralNetsweightVec_40),
    .io_out_bits_confneuralNetsweightVec_41(configurationMemory_io_out_bits_confneuralNetsweightVec_41),
    .io_out_bits_confneuralNetsweightVec_42(configurationMemory_io_out_bits_confneuralNetsweightVec_42),
    .io_out_bits_confneuralNetsweightVec_43(configurationMemory_io_out_bits_confneuralNetsweightVec_43),
    .io_out_bits_confneuralNetsweightVec_44(configurationMemory_io_out_bits_confneuralNetsweightVec_44),
    .io_out_bits_confneuralNetsweightVec_45(configurationMemory_io_out_bits_confneuralNetsweightVec_45),
    .io_out_bits_confneuralNetsweightVec_46(configurationMemory_io_out_bits_confneuralNetsweightVec_46),
    .io_out_bits_confneuralNetsweightVec_47(configurationMemory_io_out_bits_confneuralNetsweightVec_47),
    .io_out_bits_confneuralNetsweightVec_48(configurationMemory_io_out_bits_confneuralNetsweightVec_48),
    .io_out_bits_confneuralNetsweightVec_49(configurationMemory_io_out_bits_confneuralNetsweightVec_49),
    .io_out_bits_confneuralNetsweightVec_50(configurationMemory_io_out_bits_confneuralNetsweightVec_50),
    .io_out_bits_confneuralNetsweightVec_51(configurationMemory_io_out_bits_confneuralNetsweightVec_51),
    .io_out_bits_confneuralNetsweightVec_52(configurationMemory_io_out_bits_confneuralNetsweightVec_52),
    .io_out_bits_confneuralNetsweightVec_53(configurationMemory_io_out_bits_confneuralNetsweightVec_53),
    .io_out_bits_confneuralNetsweightVec_54(configurationMemory_io_out_bits_confneuralNetsweightVec_54),
    .io_out_bits_confneuralNetsweightVec_55(configurationMemory_io_out_bits_confneuralNetsweightVec_55),
    .io_out_bits_confneuralNetsweightVec_56(configurationMemory_io_out_bits_confneuralNetsweightVec_56),
    .io_out_bits_confneuralNetsweightVec_57(configurationMemory_io_out_bits_confneuralNetsweightVec_57),
    .io_out_bits_confneuralNetsweightVec_58(configurationMemory_io_out_bits_confneuralNetsweightVec_58),
    .io_out_bits_confneuralNetsweightVec_59(configurationMemory_io_out_bits_confneuralNetsweightVec_59),
    .io_out_bits_confneuralNetsweightVec_60(configurationMemory_io_out_bits_confneuralNetsweightVec_60),
    .io_out_bits_confneuralNetsweightVec_61(configurationMemory_io_out_bits_confneuralNetsweightVec_61),
    .io_out_bits_confneuralNetsweightVec_62(configurationMemory_io_out_bits_confneuralNetsweightVec_62),
    .io_out_bits_confneuralNetsweightVec_63(configurationMemory_io_out_bits_confneuralNetsweightVec_63),
    .io_out_bits_confneuralNetsweightVec_64(configurationMemory_io_out_bits_confneuralNetsweightVec_64),
    .io_out_bits_confneuralNetsweightVec_65(configurationMemory_io_out_bits_confneuralNetsweightVec_65),
    .io_out_bits_confneuralNetsweightVec_66(configurationMemory_io_out_bits_confneuralNetsweightVec_66),
    .io_out_bits_confneuralNetsweightVec_67(configurationMemory_io_out_bits_confneuralNetsweightVec_67),
    .io_out_bits_confneuralNetsweightVec_68(configurationMemory_io_out_bits_confneuralNetsweightVec_68),
    .io_out_bits_confneuralNetsweightVec_69(configurationMemory_io_out_bits_confneuralNetsweightVec_69),
    .io_out_bits_confneuralNetsweightVec_70(configurationMemory_io_out_bits_confneuralNetsweightVec_70),
    .io_out_bits_confneuralNetsweightVec_71(configurationMemory_io_out_bits_confneuralNetsweightVec_71),
    .io_out_bits_confneuralNetsweightVec_72(configurationMemory_io_out_bits_confneuralNetsweightVec_72),
    .io_out_bits_confneuralNetsweightVec_73(configurationMemory_io_out_bits_confneuralNetsweightVec_73),
    .io_out_bits_confneuralNetsweightVec_74(configurationMemory_io_out_bits_confneuralNetsweightVec_74),
    .io_out_bits_confneuralNetsweightVec_75(configurationMemory_io_out_bits_confneuralNetsweightVec_75),
    .io_out_bits_confneuralNetsweightVec_76(configurationMemory_io_out_bits_confneuralNetsweightVec_76),
    .io_out_bits_confneuralNetsweightVec_77(configurationMemory_io_out_bits_confneuralNetsweightVec_77),
    .io_out_bits_confneuralNetsweightVec_78(configurationMemory_io_out_bits_confneuralNetsweightVec_78),
    .io_out_bits_confneuralNetsweightVec_79(configurationMemory_io_out_bits_confneuralNetsweightVec_79),
    .io_out_bits_confneuralNetsweightVec_80(configurationMemory_io_out_bits_confneuralNetsweightVec_80),
    .io_out_bits_confneuralNetsweightVec_81(configurationMemory_io_out_bits_confneuralNetsweightVec_81),
    .io_out_bits_confneuralNetsweightVec_82(configurationMemory_io_out_bits_confneuralNetsweightVec_82),
    .io_out_bits_confneuralNetsweightVec_83(configurationMemory_io_out_bits_confneuralNetsweightVec_83),
    .io_out_bits_confneuralNetsweightVec_84(configurationMemory_io_out_bits_confneuralNetsweightVec_84),
    .io_out_bits_confneuralNetsweightVec_85(configurationMemory_io_out_bits_confneuralNetsweightVec_85),
    .io_out_bits_confneuralNetsweightVec_86(configurationMemory_io_out_bits_confneuralNetsweightVec_86),
    .io_out_bits_confneuralNetsweightVec_87(configurationMemory_io_out_bits_confneuralNetsweightVec_87),
    .io_out_bits_confneuralNetsweightVec_88(configurationMemory_io_out_bits_confneuralNetsweightVec_88),
    .io_out_bits_confneuralNetsweightVec_89(configurationMemory_io_out_bits_confneuralNetsweightVec_89),
    .io_out_bits_confneuralNetsweightVec_90(configurationMemory_io_out_bits_confneuralNetsweightVec_90),
    .io_out_bits_confneuralNetsweightVec_91(configurationMemory_io_out_bits_confneuralNetsweightVec_91),
    .io_out_bits_confneuralNetsweightVec_92(configurationMemory_io_out_bits_confneuralNetsweightVec_92),
    .io_out_bits_confneuralNetsweightVec_93(configurationMemory_io_out_bits_confneuralNetsweightVec_93),
    .io_out_bits_confneuralNetsweightVec_94(configurationMemory_io_out_bits_confneuralNetsweightVec_94),
    .io_out_bits_confneuralNetsweightVec_95(configurationMemory_io_out_bits_confneuralNetsweightVec_95),
    .io_out_bits_confneuralNetsweightVec_96(configurationMemory_io_out_bits_confneuralNetsweightVec_96),
    .io_out_bits_confneuralNetsweightVec_97(configurationMemory_io_out_bits_confneuralNetsweightVec_97),
    .io_out_bits_confneuralNetsweightVec_98(configurationMemory_io_out_bits_confneuralNetsweightVec_98),
    .io_out_bits_confneuralNetsweightVec_99(configurationMemory_io_out_bits_confneuralNetsweightVec_99),
    .io_out_bits_confneuralNetsbiasVec_0(configurationMemory_io_out_bits_confneuralNetsbiasVec_0),
    .io_out_bits_confneuralNetsbiasVec_1(configurationMemory_io_out_bits_confneuralNetsbiasVec_1),
    .io_out_bits_confneuralNetsbiasVec_2(configurationMemory_io_out_bits_confneuralNetsbiasVec_2),
    .io_out_bits_confneuralNetsbiasVec_3(configurationMemory_io_out_bits_confneuralNetsbiasVec_3),
    .io_out_bits_confneuralNetsbiasVec_4(configurationMemory_io_out_bits_confneuralNetsbiasVec_4),
    .io_out_bits_confneuralNetsbiasVec_5(configurationMemory_io_out_bits_confneuralNetsbiasVec_5),
    .io_out_bits_confneuralNetsbiasVec_6(configurationMemory_io_out_bits_confneuralNetsbiasVec_6),
    .io_out_bits_confneuralNetsbiasVec_7(configurationMemory_io_out_bits_confneuralNetsbiasVec_7),
    .io_out_bits_confneuralNetsbiasVec_8(configurationMemory_io_out_bits_confneuralNetsbiasVec_8),
    .io_out_bits_confneuralNetsbiasVec_9(configurationMemory_io_out_bits_confneuralNetsbiasVec_9),
    .io_out_bits_confneuralNetsbiasVec_10(configurationMemory_io_out_bits_confneuralNetsbiasVec_10),
    .io_out_bits_confneuralNetsbiasVec_11(configurationMemory_io_out_bits_confneuralNetsbiasVec_11),
    .io_out_bits_confneuralNetsbiasVec_12(configurationMemory_io_out_bits_confneuralNetsbiasVec_12),
    .io_out_bits_confneuralNetsbiasVec_13(configurationMemory_io_out_bits_confneuralNetsbiasVec_13),
    .io_out_bits_confneuralNetsbiasVec_14(configurationMemory_io_out_bits_confneuralNetsbiasVec_14),
    .io_out_bits_confneuralNetsbiasVec_15(configurationMemory_io_out_bits_confneuralNetsbiasVec_15),
    .io_out_bits_confneuralNetsbiasVec_16(configurationMemory_io_out_bits_confneuralNetsbiasVec_16),
    .io_out_bits_confneuralNetsbiasVec_17(configurationMemory_io_out_bits_confneuralNetsbiasVec_17),
    .io_out_bits_confneuralNetsbiasVec_18(configurationMemory_io_out_bits_confneuralNetsbiasVec_18),
    .io_out_bits_confneuralNetsbiasVec_19(configurationMemory_io_out_bits_confneuralNetsbiasVec_19),
    .io_out_bits_confneuralNetsbiasVec_20(configurationMemory_io_out_bits_confneuralNetsbiasVec_20),
    .io_out_bits_confneuralNetsbiasVec_21(configurationMemory_io_out_bits_confneuralNetsbiasVec_21),
    .io_out_bits_confneuralNetsbiasVec_22(configurationMemory_io_out_bits_confneuralNetsbiasVec_22),
    .io_out_bits_confneuralNetsbiasVec_23(configurationMemory_io_out_bits_confneuralNetsbiasVec_23),
    .io_out_bits_confneuralNetsbiasVec_24(configurationMemory_io_out_bits_confneuralNetsbiasVec_24),
    .io_out_bits_confneuralNetsbiasVec_25(configurationMemory_io_out_bits_confneuralNetsbiasVec_25),
    .io_out_bits_confneuralNetsbiasVec_26(configurationMemory_io_out_bits_confneuralNetsbiasVec_26),
    .io_out_bits_confneuralNetsbiasVec_27(configurationMemory_io_out_bits_confneuralNetsbiasVec_27),
    .io_out_bits_confneuralNetsbiasVec_28(configurationMemory_io_out_bits_confneuralNetsbiasVec_28),
    .io_out_bits_confneuralNetsbiasVec_29(configurationMemory_io_out_bits_confneuralNetsbiasVec_29),
    .io_out_bits_confneuralNetsbiasVec_30(configurationMemory_io_out_bits_confneuralNetsbiasVec_30),
    .io_out_bits_confneuralNetsbiasVec_31(configurationMemory_io_out_bits_confneuralNetsbiasVec_31),
    .io_out_bits_confneuralNetsbiasVec_32(configurationMemory_io_out_bits_confneuralNetsbiasVec_32),
    .io_out_bits_confneuralNetsbiasVec_33(configurationMemory_io_out_bits_confneuralNetsbiasVec_33),
    .io_out_bits_confneuralNetsbiasVec_34(configurationMemory_io_out_bits_confneuralNetsbiasVec_34),
    .io_out_bits_confneuralNetsbiasVec_35(configurationMemory_io_out_bits_confneuralNetsbiasVec_35),
    .io_out_bits_confneuralNetsbiasVec_36(configurationMemory_io_out_bits_confneuralNetsbiasVec_36),
    .io_out_bits_confneuralNetsbiasVec_37(configurationMemory_io_out_bits_confneuralNetsbiasVec_37),
    .io_out_bits_confneuralNetsbiasVec_38(configurationMemory_io_out_bits_confneuralNetsbiasVec_38),
    .io_out_bits_confneuralNetsbiasVec_39(configurationMemory_io_out_bits_confneuralNetsbiasVec_39),
    .io_out_bits_confneuralNetsbiasVec_40(configurationMemory_io_out_bits_confneuralNetsbiasVec_40),
    .io_out_bits_confneuralNetsbiasVec_41(configurationMemory_io_out_bits_confneuralNetsbiasVec_41),
    .io_out_bits_confneuralNetsbiasVec_42(configurationMemory_io_out_bits_confneuralNetsbiasVec_42),
    .io_out_bits_confneuralNetsbiasVec_43(configurationMemory_io_out_bits_confneuralNetsbiasVec_43),
    .io_out_bits_confneuralNetsbiasVec_44(configurationMemory_io_out_bits_confneuralNetsbiasVec_44),
    .io_out_bits_confneuralNetsbiasVec_45(configurationMemory_io_out_bits_confneuralNetsbiasVec_45),
    .io_out_bits_confneuralNetsbiasVec_46(configurationMemory_io_out_bits_confneuralNetsbiasVec_46),
    .io_out_bits_confneuralNetsbiasVec_47(configurationMemory_io_out_bits_confneuralNetsbiasVec_47),
    .io_out_bits_confneuralNetsbiasVec_48(configurationMemory_io_out_bits_confneuralNetsbiasVec_48),
    .io_out_bits_confneuralNetsbiasVec_49(configurationMemory_io_out_bits_confneuralNetsbiasVec_49),
    .io_out_bits_confneuralNetsbiasVec_50(configurationMemory_io_out_bits_confneuralNetsbiasVec_50),
    .io_out_bits_confneuralNetsbiasVec_51(configurationMemory_io_out_bits_confneuralNetsbiasVec_51),
    .io_out_bits_confneuralNetsbiasVec_52(configurationMemory_io_out_bits_confneuralNetsbiasVec_52),
    .io_out_bits_confneuralNetsbiasVec_53(configurationMemory_io_out_bits_confneuralNetsbiasVec_53),
    .io_out_bits_confneuralNetsbiasVec_54(configurationMemory_io_out_bits_confneuralNetsbiasVec_54),
    .io_out_bits_confneuralNetsbiasVec_55(configurationMemory_io_out_bits_confneuralNetsbiasVec_55),
    .io_out_bits_confneuralNetsbiasVec_56(configurationMemory_io_out_bits_confneuralNetsbiasVec_56),
    .io_out_bits_confneuralNetsbiasVec_57(configurationMemory_io_out_bits_confneuralNetsbiasVec_57),
    .io_out_bits_confneuralNetsbiasVec_58(configurationMemory_io_out_bits_confneuralNetsbiasVec_58),
    .io_out_bits_confneuralNetsbiasVec_59(configurationMemory_io_out_bits_confneuralNetsbiasVec_59),
    .io_out_bits_confneuralNetsbiasVec_60(configurationMemory_io_out_bits_confneuralNetsbiasVec_60),
    .io_out_bits_confneuralNetsbiasVec_61(configurationMemory_io_out_bits_confneuralNetsbiasVec_61),
    .io_out_bits_confneuralNetsbiasVec_62(configurationMemory_io_out_bits_confneuralNetsbiasVec_62),
    .io_out_bits_confneuralNetsbiasVec_63(configurationMemory_io_out_bits_confneuralNetsbiasVec_63),
    .io_out_bits_confneuralNetsbiasVec_64(configurationMemory_io_out_bits_confneuralNetsbiasVec_64),
    .io_out_bits_confneuralNetsbiasVec_65(configurationMemory_io_out_bits_confneuralNetsbiasVec_65),
    .io_out_bits_confneuralNetsbiasVec_66(configurationMemory_io_out_bits_confneuralNetsbiasVec_66),
    .io_out_bits_confneuralNetsbiasVec_67(configurationMemory_io_out_bits_confneuralNetsbiasVec_67),
    .io_out_bits_confneuralNetsbiasVec_68(configurationMemory_io_out_bits_confneuralNetsbiasVec_68),
    .io_out_bits_confneuralNetsbiasVec_69(configurationMemory_io_out_bits_confneuralNetsbiasVec_69),
    .io_out_bits_confneuralNetsbiasVec_70(configurationMemory_io_out_bits_confneuralNetsbiasVec_70),
    .io_out_bits_confneuralNetsbiasVec_71(configurationMemory_io_out_bits_confneuralNetsbiasVec_71),
    .io_out_bits_confneuralNetsbiasVec_72(configurationMemory_io_out_bits_confneuralNetsbiasVec_72),
    .io_out_bits_confneuralNetsbiasVec_73(configurationMemory_io_out_bits_confneuralNetsbiasVec_73),
    .io_out_bits_confneuralNetsbiasVec_74(configurationMemory_io_out_bits_confneuralNetsbiasVec_74),
    .io_out_bits_confneuralNetsbiasVec_75(configurationMemory_io_out_bits_confneuralNetsbiasVec_75),
    .io_out_bits_confneuralNetsbiasVec_76(configurationMemory_io_out_bits_confneuralNetsbiasVec_76),
    .io_out_bits_confneuralNetsbiasVec_77(configurationMemory_io_out_bits_confneuralNetsbiasVec_77),
    .io_out_bits_confneuralNetsbiasVec_78(configurationMemory_io_out_bits_confneuralNetsbiasVec_78),
    .io_out_bits_confneuralNetsbiasVec_79(configurationMemory_io_out_bits_confneuralNetsbiasVec_79),
    .io_out_bits_confneuralNetsbiasVec_80(configurationMemory_io_out_bits_confneuralNetsbiasVec_80),
    .io_out_bits_confneuralNetsbiasVec_81(configurationMemory_io_out_bits_confneuralNetsbiasVec_81),
    .io_out_bits_confneuralNetsbiasVec_82(configurationMemory_io_out_bits_confneuralNetsbiasVec_82),
    .io_out_bits_confneuralNetsbiasVec_83(configurationMemory_io_out_bits_confneuralNetsbiasVec_83),
    .io_out_bits_confneuralNetsbiasVec_84(configurationMemory_io_out_bits_confneuralNetsbiasVec_84),
    .io_out_bits_confneuralNetsbiasVec_85(configurationMemory_io_out_bits_confneuralNetsbiasVec_85),
    .io_out_bits_confneuralNetsbiasVec_86(configurationMemory_io_out_bits_confneuralNetsbiasVec_86),
    .io_out_bits_confneuralNetsbiasVec_87(configurationMemory_io_out_bits_confneuralNetsbiasVec_87),
    .io_out_bits_confneuralNetsbiasVec_88(configurationMemory_io_out_bits_confneuralNetsbiasVec_88),
    .io_out_bits_confneuralNetsbiasVec_89(configurationMemory_io_out_bits_confneuralNetsbiasVec_89),
    .io_out_bits_confneuralNetsbiasVec_90(configurationMemory_io_out_bits_confneuralNetsbiasVec_90),
    .io_out_bits_confneuralNetsbiasVec_91(configurationMemory_io_out_bits_confneuralNetsbiasVec_91),
    .io_out_bits_confneuralNetsbiasVec_92(configurationMemory_io_out_bits_confneuralNetsbiasVec_92),
    .io_out_bits_confneuralNetsbiasVec_93(configurationMemory_io_out_bits_confneuralNetsbiasVec_93),
    .io_out_bits_confneuralNetsbiasVec_94(configurationMemory_io_out_bits_confneuralNetsbiasVec_94),
    .io_out_bits_confneuralNetsbiasVec_95(configurationMemory_io_out_bits_confneuralNetsbiasVec_95),
    .io_out_bits_confneuralNetsbiasVec_96(configurationMemory_io_out_bits_confneuralNetsbiasVec_96),
    .io_out_bits_confneuralNetsbiasVec_97(configurationMemory_io_out_bits_confneuralNetsbiasVec_97),
    .io_out_bits_confneuralNetsbiasVec_98(configurationMemory_io_out_bits_confneuralNetsbiasVec_98),
    .io_out_bits_confneuralNetsbiasVec_99(configurationMemory_io_out_bits_confneuralNetsbiasVec_99),
    .io_out_bits_confneuralNetsbiasScalar_0(configurationMemory_io_out_bits_confneuralNetsbiasScalar_0),
    .io_out_bits_confInputMuxSel(configurationMemory_io_out_bits_confInputMuxSel)
  );
  assign in_1_bits_data = converter_1_auto_out_bits_data; // @[Nodes.scala 333:76 LazyModule.scala 167:31]
  assign _T_4 = $signed(in_1_bits_data); // @[Wellness.scala 408:49]
  assign _T_5 = $unsigned(wellness_io_rawVotes); // @[Wellness.scala 411:83]
  assign _T_6 = {wellness_io_out_bits,_T_5}; // @[Cat.scala 30:58]
  assign inConf_bits_data = converter_2_auto_out_bits_data; // @[Nodes.scala 333:76 LazyModule.scala 167:31]
  assign _T_7 = inConf_bits_data[31:0]; // @[Wellness.scala 418:62]
  assign _GEN_0 = _T_4[31:0]; // @[Wellness.scala 408:49 Wellness.scala 408:49]
  assign in_ready = converter_1_auto_in_ready; // @[BundleBridge.scala 39:12]
  assign out_valid = converter_auto_out_valid; // @[BundleBridge.scala 27:8]
  assign out_bits_data = converter_auto_out_bits_data; // @[BundleBridge.scala 27:8]
  assign out_bits_last = converter_auto_out_bits_last; // @[BundleBridge.scala 27:8]
  assign in2_ready = converter_2_auto_in_ready; // @[BundleBridge.scala 39:12]
  assign converter_auto_in_valid = wellness_io_out_valid; // @[LazyModule.scala 167:57]
  assign converter_auto_in_bits_data = {{31'd0}, _T_6}; // @[LazyModule.scala 167:57]
  assign converter_auto_in_bits_last = 1'h0; // @[LazyModule.scala 167:57]
  assign converter_auto_out_ready = out_ready; // @[LazyModule.scala 167:31]
  assign converter_1_auto_in_valid = in_valid; // @[LazyModule.scala 167:57]
  assign converter_1_auto_in_bits_data = in_bits_data; // @[LazyModule.scala 167:57]
  assign converter_1_auto_in_bits_last = in_bits_last; // @[LazyModule.scala 167:57]
  assign converter_1_auto_out_ready = 1'h1; // @[LazyModule.scala 167:31]
  assign converter_2_auto_in_valid = in2_valid; // @[LazyModule.scala 167:57]
  assign converter_2_auto_in_bits_data = in2_bits_data; // @[LazyModule.scala 167:57]
  assign converter_2_auto_in_bits_last = in2_bits_last; // @[LazyModule.scala 167:57]
  assign converter_2_auto_out_ready = 1'h1; // @[LazyModule.scala 167:31]
  assign wellness_clock = clock;
  assign wellness_reset = reset;
  assign wellness_io_streamIn_valid = streamIn_valid; // @[Wellness.scala 402:32]
  assign wellness_io_streamIn_bits = streamIn_bits; // @[Wellness.scala 401:31]
  assign wellness_io_in_valid = converter_1_auto_out_valid; // @[Wellness.scala 407:26]
  assign wellness_io_in_bits = $signed(_GEN_0); // @[Wellness.scala 408:25]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_0_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_0_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_0_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_0_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_0_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_0_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_0_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_0_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_1_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_1_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_1_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_1_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_1_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_1_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_1_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_1_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_2_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_2_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_2_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_2_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_2_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_2_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_2_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_2_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_3_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_3_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_3_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_3_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_3_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_3_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_3_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_3_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_4_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_4_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_4_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_4_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_4_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_4_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_4_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_4_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_5_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_5_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_5_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_5_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_5_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_5_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_5_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_5_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_6_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_6_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_6_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_6_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_6_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_6_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_6_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_6_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_7_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_7_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_7_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_7_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_7_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_7_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_7_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_7_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_8_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_8_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_8_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_8_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_8_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_8_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_8_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_8_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_9_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_9_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_9_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_9_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_9_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_9_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_9_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_9_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_10_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_10_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_10_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_10_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_10_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_10_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_10_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_10_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_11_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_11_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_11_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_11_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_11_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_11_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_11_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_11_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_12_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_12_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_12_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_12_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_12_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_12_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_12_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_12_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_13_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_13_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_13_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_13_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_13_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_13_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_13_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_13_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_14_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_14_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_14_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_14_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_14_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_14_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_14_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_14_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_15_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_15_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_15_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_15_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_15_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_15_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_15_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_15_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_16_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_16_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_16_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_16_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_16_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_16_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_16_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_16_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_17_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_17_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_17_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_17_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_17_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_17_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_17_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_17_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_18_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_18_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_18_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_18_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_18_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_18_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_18_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_18_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_19_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_19_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_19_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_19_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_19_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_19_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_19_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_19_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_20_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_20_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_20_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_20_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_20_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_20_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_20_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_20_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_21_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_21_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_21_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_21_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_21_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_21_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_21_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_21_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_22_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_22_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_22_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_22_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_22_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_22_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_22_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_22_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_23_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_23_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_23_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_23_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_23_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_23_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_23_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_23_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_24_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_24_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_24_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_24_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_24_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_24_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_24_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_24_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_25_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_25_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_25_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_25_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_25_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_25_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_25_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_25_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_26_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_26_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_26_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_26_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_26_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_26_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_26_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_26_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_27_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_27_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_27_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_27_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_27_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_27_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_27_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_27_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_28_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_28_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_28_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_28_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_28_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_28_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_28_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_28_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_29_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_29_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_29_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_29_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_29_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_29_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_29_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_29_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_30_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_30_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_30_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_30_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_30_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_30_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_30_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_30_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_31_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_31_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_31_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_31_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_31_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_31_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_31_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_31_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_32_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_32_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_32_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_32_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_32_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_32_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_32_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_32_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_33_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_33_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_33_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_33_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_33_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_33_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_33_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_33_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_34_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_34_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_34_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_34_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_34_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_34_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_34_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_34_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_35_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_35_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_35_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_35_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_35_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_35_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_35_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_35_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_36_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_36_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_36_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_36_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_36_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_36_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_36_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_36_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_37_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_37_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_37_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_37_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_37_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_37_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_37_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_37_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_38_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_38_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_38_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_38_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_38_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_38_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_38_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_38_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_39_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_39_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_39_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_39_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_39_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_39_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_39_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_39_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_40_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_40_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_40_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_40_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_40_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_40_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_40_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_40_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_41_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_41_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_41_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_41_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_41_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_41_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_41_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_41_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_42_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_42_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_42_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_42_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_42_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_42_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_42_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_42_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_43_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_43_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_43_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_43_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_43_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_43_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_43_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_43_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_44_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_44_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_44_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_44_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_44_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_44_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_44_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_44_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_45_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_45_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_45_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_45_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_45_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_45_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_45_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_45_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_46_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_46_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_46_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_46_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_46_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_46_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_46_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_46_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_47_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_47_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_47_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_47_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_47_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_47_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_47_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_47_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_48_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_48_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_48_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_48_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_48_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_48_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_48_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_48_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_49_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_49_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_49_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_49_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_49_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_49_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_49_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_49_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_50_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_50_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_50_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_50_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_50_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_50_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_50_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_50_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_51_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_51_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_51_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_51_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_51_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_51_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_51_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_51_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_52_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_52_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_52_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_52_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_52_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_52_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_52_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_52_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_53_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_53_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_53_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_53_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_53_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_53_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_53_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_53_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_54_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_54_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_54_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_54_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_54_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_54_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_54_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_54_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_55_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_55_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_55_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_55_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_55_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_55_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_55_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_55_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_56_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_56_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_56_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_56_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_56_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_56_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_56_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_56_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_57_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_57_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_57_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_57_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_57_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_57_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_57_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_57_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_58_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_58_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_58_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_58_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_58_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_58_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_58_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_58_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_59_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_59_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_59_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_59_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_59_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_59_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_59_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_59_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_60_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_60_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_60_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_60_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_60_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_60_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_60_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_60_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_61_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_61_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_61_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_61_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_61_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_61_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_61_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_61_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_62_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_62_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_62_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_62_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_62_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_62_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_62_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_62_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_63_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_63_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_63_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_63_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_63_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_63_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_63_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_63_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_64_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_64_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_64_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_64_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_64_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_64_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_64_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_64_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_65_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_65_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_65_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_65_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_65_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_65_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_65_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_65_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_66_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_66_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_66_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_66_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_66_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_66_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_66_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_66_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_67_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_67_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_67_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_67_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_67_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_67_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_67_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_67_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_68_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_68_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_68_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_68_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_68_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_68_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_68_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_68_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_69_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_69_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_69_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_69_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_69_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_69_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_69_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_69_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_70_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_70_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_70_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_70_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_70_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_70_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_70_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_70_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_71_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_71_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_71_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_71_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_71_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_71_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_71_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_71_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_72_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_72_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_72_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_72_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_72_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_72_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_72_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_72_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_73_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_73_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_73_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_73_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_73_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_73_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_73_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_73_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_74_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_74_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_74_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_74_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_74_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_74_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_74_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_74_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_75_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_75_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_75_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_75_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_75_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_75_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_75_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_75_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_76_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_76_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_76_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_76_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_76_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_76_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_76_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_76_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_77_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_77_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_77_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_77_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_77_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_77_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_77_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_77_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_78_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_78_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_78_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_78_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_78_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_78_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_78_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_78_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_79_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_79_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_79_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_79_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_79_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_79_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_79_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_79_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_80_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_80_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_80_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_80_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_80_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_80_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_80_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_80_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_81_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_81_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_81_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_81_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_81_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_81_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_81_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_81_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_82_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_82_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_82_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_82_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_82_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_82_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_82_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_82_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_83_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_83_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_83_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_83_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_83_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_83_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_83_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_83_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_84_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_84_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_84_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_84_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_84_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_84_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_84_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_84_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_85_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_85_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_85_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_85_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_85_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_85_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_85_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_85_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_86_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_86_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_86_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_86_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_86_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_86_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_86_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_86_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_87_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_87_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_87_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_87_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_87_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_87_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_87_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_87_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_88_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_88_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_88_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_88_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_88_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_88_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_88_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_88_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_89_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_89_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_89_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_89_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_89_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_89_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_89_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_89_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_90_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_90_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_90_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_90_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_90_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_90_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_90_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_90_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_91_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_91_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_91_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_91_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_91_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_91_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_91_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_91_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_92_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_92_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_92_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_92_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_92_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_92_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_92_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_92_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_93_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_93_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_93_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_93_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_93_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_93_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_93_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_93_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_94_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_94_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_94_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_94_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_94_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_94_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_94_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_94_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_95_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_95_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_95_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_95_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_95_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_95_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_95_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_95_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_96_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_96_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_96_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_96_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_96_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_96_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_96_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_96_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_97_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_97_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_97_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_97_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_97_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_97_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_97_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_97_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_98_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_98_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_98_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_98_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_98_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_98_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_98_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_98_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_99_0 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_99_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_99_1 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_99_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_99_2 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_99_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightMatrix_99_3 = configurationMemory_io_out_bits_confneuralNetsweightMatrix_99_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_0 = configurationMemory_io_out_bits_confneuralNetsweightVec_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_1 = configurationMemory_io_out_bits_confneuralNetsweightVec_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_2 = configurationMemory_io_out_bits_confneuralNetsweightVec_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_3 = configurationMemory_io_out_bits_confneuralNetsweightVec_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_4 = configurationMemory_io_out_bits_confneuralNetsweightVec_4; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_5 = configurationMemory_io_out_bits_confneuralNetsweightVec_5; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_6 = configurationMemory_io_out_bits_confneuralNetsweightVec_6; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_7 = configurationMemory_io_out_bits_confneuralNetsweightVec_7; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_8 = configurationMemory_io_out_bits_confneuralNetsweightVec_8; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_9 = configurationMemory_io_out_bits_confneuralNetsweightVec_9; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_10 = configurationMemory_io_out_bits_confneuralNetsweightVec_10; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_11 = configurationMemory_io_out_bits_confneuralNetsweightVec_11; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_12 = configurationMemory_io_out_bits_confneuralNetsweightVec_12; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_13 = configurationMemory_io_out_bits_confneuralNetsweightVec_13; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_14 = configurationMemory_io_out_bits_confneuralNetsweightVec_14; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_15 = configurationMemory_io_out_bits_confneuralNetsweightVec_15; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_16 = configurationMemory_io_out_bits_confneuralNetsweightVec_16; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_17 = configurationMemory_io_out_bits_confneuralNetsweightVec_17; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_18 = configurationMemory_io_out_bits_confneuralNetsweightVec_18; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_19 = configurationMemory_io_out_bits_confneuralNetsweightVec_19; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_20 = configurationMemory_io_out_bits_confneuralNetsweightVec_20; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_21 = configurationMemory_io_out_bits_confneuralNetsweightVec_21; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_22 = configurationMemory_io_out_bits_confneuralNetsweightVec_22; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_23 = configurationMemory_io_out_bits_confneuralNetsweightVec_23; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_24 = configurationMemory_io_out_bits_confneuralNetsweightVec_24; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_25 = configurationMemory_io_out_bits_confneuralNetsweightVec_25; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_26 = configurationMemory_io_out_bits_confneuralNetsweightVec_26; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_27 = configurationMemory_io_out_bits_confneuralNetsweightVec_27; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_28 = configurationMemory_io_out_bits_confneuralNetsweightVec_28; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_29 = configurationMemory_io_out_bits_confneuralNetsweightVec_29; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_30 = configurationMemory_io_out_bits_confneuralNetsweightVec_30; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_31 = configurationMemory_io_out_bits_confneuralNetsweightVec_31; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_32 = configurationMemory_io_out_bits_confneuralNetsweightVec_32; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_33 = configurationMemory_io_out_bits_confneuralNetsweightVec_33; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_34 = configurationMemory_io_out_bits_confneuralNetsweightVec_34; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_35 = configurationMemory_io_out_bits_confneuralNetsweightVec_35; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_36 = configurationMemory_io_out_bits_confneuralNetsweightVec_36; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_37 = configurationMemory_io_out_bits_confneuralNetsweightVec_37; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_38 = configurationMemory_io_out_bits_confneuralNetsweightVec_38; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_39 = configurationMemory_io_out_bits_confneuralNetsweightVec_39; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_40 = configurationMemory_io_out_bits_confneuralNetsweightVec_40; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_41 = configurationMemory_io_out_bits_confneuralNetsweightVec_41; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_42 = configurationMemory_io_out_bits_confneuralNetsweightVec_42; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_43 = configurationMemory_io_out_bits_confneuralNetsweightVec_43; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_44 = configurationMemory_io_out_bits_confneuralNetsweightVec_44; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_45 = configurationMemory_io_out_bits_confneuralNetsweightVec_45; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_46 = configurationMemory_io_out_bits_confneuralNetsweightVec_46; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_47 = configurationMemory_io_out_bits_confneuralNetsweightVec_47; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_48 = configurationMemory_io_out_bits_confneuralNetsweightVec_48; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_49 = configurationMemory_io_out_bits_confneuralNetsweightVec_49; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_50 = configurationMemory_io_out_bits_confneuralNetsweightVec_50; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_51 = configurationMemory_io_out_bits_confneuralNetsweightVec_51; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_52 = configurationMemory_io_out_bits_confneuralNetsweightVec_52; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_53 = configurationMemory_io_out_bits_confneuralNetsweightVec_53; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_54 = configurationMemory_io_out_bits_confneuralNetsweightVec_54; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_55 = configurationMemory_io_out_bits_confneuralNetsweightVec_55; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_56 = configurationMemory_io_out_bits_confneuralNetsweightVec_56; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_57 = configurationMemory_io_out_bits_confneuralNetsweightVec_57; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_58 = configurationMemory_io_out_bits_confneuralNetsweightVec_58; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_59 = configurationMemory_io_out_bits_confneuralNetsweightVec_59; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_60 = configurationMemory_io_out_bits_confneuralNetsweightVec_60; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_61 = configurationMemory_io_out_bits_confneuralNetsweightVec_61; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_62 = configurationMemory_io_out_bits_confneuralNetsweightVec_62; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_63 = configurationMemory_io_out_bits_confneuralNetsweightVec_63; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_64 = configurationMemory_io_out_bits_confneuralNetsweightVec_64; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_65 = configurationMemory_io_out_bits_confneuralNetsweightVec_65; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_66 = configurationMemory_io_out_bits_confneuralNetsweightVec_66; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_67 = configurationMemory_io_out_bits_confneuralNetsweightVec_67; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_68 = configurationMemory_io_out_bits_confneuralNetsweightVec_68; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_69 = configurationMemory_io_out_bits_confneuralNetsweightVec_69; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_70 = configurationMemory_io_out_bits_confneuralNetsweightVec_70; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_71 = configurationMemory_io_out_bits_confneuralNetsweightVec_71; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_72 = configurationMemory_io_out_bits_confneuralNetsweightVec_72; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_73 = configurationMemory_io_out_bits_confneuralNetsweightVec_73; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_74 = configurationMemory_io_out_bits_confneuralNetsweightVec_74; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_75 = configurationMemory_io_out_bits_confneuralNetsweightVec_75; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_76 = configurationMemory_io_out_bits_confneuralNetsweightVec_76; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_77 = configurationMemory_io_out_bits_confneuralNetsweightVec_77; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_78 = configurationMemory_io_out_bits_confneuralNetsweightVec_78; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_79 = configurationMemory_io_out_bits_confneuralNetsweightVec_79; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_80 = configurationMemory_io_out_bits_confneuralNetsweightVec_80; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_81 = configurationMemory_io_out_bits_confneuralNetsweightVec_81; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_82 = configurationMemory_io_out_bits_confneuralNetsweightVec_82; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_83 = configurationMemory_io_out_bits_confneuralNetsweightVec_83; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_84 = configurationMemory_io_out_bits_confneuralNetsweightVec_84; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_85 = configurationMemory_io_out_bits_confneuralNetsweightVec_85; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_86 = configurationMemory_io_out_bits_confneuralNetsweightVec_86; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_87 = configurationMemory_io_out_bits_confneuralNetsweightVec_87; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_88 = configurationMemory_io_out_bits_confneuralNetsweightVec_88; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_89 = configurationMemory_io_out_bits_confneuralNetsweightVec_89; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_90 = configurationMemory_io_out_bits_confneuralNetsweightVec_90; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_91 = configurationMemory_io_out_bits_confneuralNetsweightVec_91; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_92 = configurationMemory_io_out_bits_confneuralNetsweightVec_92; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_93 = configurationMemory_io_out_bits_confneuralNetsweightVec_93; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_94 = configurationMemory_io_out_bits_confneuralNetsweightVec_94; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_95 = configurationMemory_io_out_bits_confneuralNetsweightVec_95; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_96 = configurationMemory_io_out_bits_confneuralNetsweightVec_96; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_97 = configurationMemory_io_out_bits_confneuralNetsweightVec_97; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_98 = configurationMemory_io_out_bits_confneuralNetsweightVec_98; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsweightVec_99 = configurationMemory_io_out_bits_confneuralNetsweightVec_99; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_0 = configurationMemory_io_out_bits_confneuralNetsbiasVec_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_1 = configurationMemory_io_out_bits_confneuralNetsbiasVec_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_2 = configurationMemory_io_out_bits_confneuralNetsbiasVec_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_3 = configurationMemory_io_out_bits_confneuralNetsbiasVec_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_4 = configurationMemory_io_out_bits_confneuralNetsbiasVec_4; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_5 = configurationMemory_io_out_bits_confneuralNetsbiasVec_5; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_6 = configurationMemory_io_out_bits_confneuralNetsbiasVec_6; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_7 = configurationMemory_io_out_bits_confneuralNetsbiasVec_7; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_8 = configurationMemory_io_out_bits_confneuralNetsbiasVec_8; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_9 = configurationMemory_io_out_bits_confneuralNetsbiasVec_9; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_10 = configurationMemory_io_out_bits_confneuralNetsbiasVec_10; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_11 = configurationMemory_io_out_bits_confneuralNetsbiasVec_11; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_12 = configurationMemory_io_out_bits_confneuralNetsbiasVec_12; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_13 = configurationMemory_io_out_bits_confneuralNetsbiasVec_13; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_14 = configurationMemory_io_out_bits_confneuralNetsbiasVec_14; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_15 = configurationMemory_io_out_bits_confneuralNetsbiasVec_15; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_16 = configurationMemory_io_out_bits_confneuralNetsbiasVec_16; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_17 = configurationMemory_io_out_bits_confneuralNetsbiasVec_17; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_18 = configurationMemory_io_out_bits_confneuralNetsbiasVec_18; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_19 = configurationMemory_io_out_bits_confneuralNetsbiasVec_19; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_20 = configurationMemory_io_out_bits_confneuralNetsbiasVec_20; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_21 = configurationMemory_io_out_bits_confneuralNetsbiasVec_21; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_22 = configurationMemory_io_out_bits_confneuralNetsbiasVec_22; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_23 = configurationMemory_io_out_bits_confneuralNetsbiasVec_23; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_24 = configurationMemory_io_out_bits_confneuralNetsbiasVec_24; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_25 = configurationMemory_io_out_bits_confneuralNetsbiasVec_25; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_26 = configurationMemory_io_out_bits_confneuralNetsbiasVec_26; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_27 = configurationMemory_io_out_bits_confneuralNetsbiasVec_27; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_28 = configurationMemory_io_out_bits_confneuralNetsbiasVec_28; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_29 = configurationMemory_io_out_bits_confneuralNetsbiasVec_29; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_30 = configurationMemory_io_out_bits_confneuralNetsbiasVec_30; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_31 = configurationMemory_io_out_bits_confneuralNetsbiasVec_31; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_32 = configurationMemory_io_out_bits_confneuralNetsbiasVec_32; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_33 = configurationMemory_io_out_bits_confneuralNetsbiasVec_33; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_34 = configurationMemory_io_out_bits_confneuralNetsbiasVec_34; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_35 = configurationMemory_io_out_bits_confneuralNetsbiasVec_35; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_36 = configurationMemory_io_out_bits_confneuralNetsbiasVec_36; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_37 = configurationMemory_io_out_bits_confneuralNetsbiasVec_37; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_38 = configurationMemory_io_out_bits_confneuralNetsbiasVec_38; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_39 = configurationMemory_io_out_bits_confneuralNetsbiasVec_39; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_40 = configurationMemory_io_out_bits_confneuralNetsbiasVec_40; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_41 = configurationMemory_io_out_bits_confneuralNetsbiasVec_41; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_42 = configurationMemory_io_out_bits_confneuralNetsbiasVec_42; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_43 = configurationMemory_io_out_bits_confneuralNetsbiasVec_43; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_44 = configurationMemory_io_out_bits_confneuralNetsbiasVec_44; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_45 = configurationMemory_io_out_bits_confneuralNetsbiasVec_45; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_46 = configurationMemory_io_out_bits_confneuralNetsbiasVec_46; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_47 = configurationMemory_io_out_bits_confneuralNetsbiasVec_47; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_48 = configurationMemory_io_out_bits_confneuralNetsbiasVec_48; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_49 = configurationMemory_io_out_bits_confneuralNetsbiasVec_49; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_50 = configurationMemory_io_out_bits_confneuralNetsbiasVec_50; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_51 = configurationMemory_io_out_bits_confneuralNetsbiasVec_51; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_52 = configurationMemory_io_out_bits_confneuralNetsbiasVec_52; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_53 = configurationMemory_io_out_bits_confneuralNetsbiasVec_53; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_54 = configurationMemory_io_out_bits_confneuralNetsbiasVec_54; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_55 = configurationMemory_io_out_bits_confneuralNetsbiasVec_55; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_56 = configurationMemory_io_out_bits_confneuralNetsbiasVec_56; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_57 = configurationMemory_io_out_bits_confneuralNetsbiasVec_57; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_58 = configurationMemory_io_out_bits_confneuralNetsbiasVec_58; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_59 = configurationMemory_io_out_bits_confneuralNetsbiasVec_59; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_60 = configurationMemory_io_out_bits_confneuralNetsbiasVec_60; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_61 = configurationMemory_io_out_bits_confneuralNetsbiasVec_61; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_62 = configurationMemory_io_out_bits_confneuralNetsbiasVec_62; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_63 = configurationMemory_io_out_bits_confneuralNetsbiasVec_63; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_64 = configurationMemory_io_out_bits_confneuralNetsbiasVec_64; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_65 = configurationMemory_io_out_bits_confneuralNetsbiasVec_65; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_66 = configurationMemory_io_out_bits_confneuralNetsbiasVec_66; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_67 = configurationMemory_io_out_bits_confneuralNetsbiasVec_67; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_68 = configurationMemory_io_out_bits_confneuralNetsbiasVec_68; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_69 = configurationMemory_io_out_bits_confneuralNetsbiasVec_69; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_70 = configurationMemory_io_out_bits_confneuralNetsbiasVec_70; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_71 = configurationMemory_io_out_bits_confneuralNetsbiasVec_71; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_72 = configurationMemory_io_out_bits_confneuralNetsbiasVec_72; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_73 = configurationMemory_io_out_bits_confneuralNetsbiasVec_73; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_74 = configurationMemory_io_out_bits_confneuralNetsbiasVec_74; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_75 = configurationMemory_io_out_bits_confneuralNetsbiasVec_75; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_76 = configurationMemory_io_out_bits_confneuralNetsbiasVec_76; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_77 = configurationMemory_io_out_bits_confneuralNetsbiasVec_77; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_78 = configurationMemory_io_out_bits_confneuralNetsbiasVec_78; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_79 = configurationMemory_io_out_bits_confneuralNetsbiasVec_79; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_80 = configurationMemory_io_out_bits_confneuralNetsbiasVec_80; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_81 = configurationMemory_io_out_bits_confneuralNetsbiasVec_81; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_82 = configurationMemory_io_out_bits_confneuralNetsbiasVec_82; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_83 = configurationMemory_io_out_bits_confneuralNetsbiasVec_83; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_84 = configurationMemory_io_out_bits_confneuralNetsbiasVec_84; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_85 = configurationMemory_io_out_bits_confneuralNetsbiasVec_85; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_86 = configurationMemory_io_out_bits_confneuralNetsbiasVec_86; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_87 = configurationMemory_io_out_bits_confneuralNetsbiasVec_87; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_88 = configurationMemory_io_out_bits_confneuralNetsbiasVec_88; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_89 = configurationMemory_io_out_bits_confneuralNetsbiasVec_89; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_90 = configurationMemory_io_out_bits_confneuralNetsbiasVec_90; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_91 = configurationMemory_io_out_bits_confneuralNetsbiasVec_91; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_92 = configurationMemory_io_out_bits_confneuralNetsbiasVec_92; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_93 = configurationMemory_io_out_bits_confneuralNetsbiasVec_93; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_94 = configurationMemory_io_out_bits_confneuralNetsbiasVec_94; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_95 = configurationMemory_io_out_bits_confneuralNetsbiasVec_95; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_96 = configurationMemory_io_out_bits_confneuralNetsbiasVec_96; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_97 = configurationMemory_io_out_bits_confneuralNetsbiasVec_97; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_98 = configurationMemory_io_out_bits_confneuralNetsbiasVec_98; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVec_99 = configurationMemory_io_out_bits_confneuralNetsbiasVec_99; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasScalar_0 = configurationMemory_io_out_bits_confneuralNetsbiasScalar_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confInputMuxSel = configurationMemory_io_out_bits_confInputMuxSel; // @[Wellness.scala 420:24]
  assign configurationMemory_clock = clock;
  assign configurationMemory_reset = reset;
  assign configurationMemory_io_in_valid = converter_2_auto_out_valid; // @[Wellness.scala 416:37]
  assign configurationMemory_io_in_bits_wrdata = $signed(_T_7); // @[Wellness.scala 418:43]
  assign configurationMemory_io_in_bits_wraddr = inConf_bits_data[34:32]; // @[Wellness.scala 419:43]
endmodule
