module AXI4StreamToBundleBridge(
  output        auto_in_ready,
  input         auto_in_valid,
  input  [63:0] auto_in_bits_data,
  input         auto_in_bits_last,
  input         auto_out_ready,
  output        auto_out_valid,
  output [63:0] auto_out_bits_data,
  output        auto_out_bits_last
);
  assign auto_in_ready = auto_out_ready; // @[LazyModule.scala 173:31]
  assign auto_out_valid = auto_in_valid; // @[LazyModule.scala 173:49]
  assign auto_out_bits_data = auto_in_bits_data; // @[LazyModule.scala 173:49]
  assign auto_out_bits_last = auto_in_bits_last; // @[LazyModule.scala 173:49]
endmodule
module ConstantCoefficientFIRFilter(
  input         clock,
  input         reset,
  input         io_in_valid,
  input  [31:0] io_in_bits,
  output        io_out_valid,
  output [31:0] io_out_bits
);
  reg [31:0] regs_0; // @[FIRFilter.scala 39:21]
  reg [31:0] _RAND_0;
  reg [31:0] regs_1; // @[FIRFilter.scala 39:21]
  reg [31:0] _RAND_1;
  reg [31:0] regs_2; // @[FIRFilter.scala 39:21]
  reg [31:0] _RAND_2;
  reg [31:0] regs_3; // @[FIRFilter.scala 39:21]
  reg [31:0] _RAND_3;
  reg [31:0] regs_4; // @[FIRFilter.scala 39:21]
  reg [31:0] _RAND_4;
  reg [31:0] regs_5; // @[FIRFilter.scala 39:21]
  reg [31:0] _RAND_5;
  wire [47:0] accumulator_0; // @[FixedPointTypeClass.scala 43:59]
  wire [48:0] muls_1; // @[FixedPointTypeClass.scala 43:59]
  wire [48:0] muls_2; // @[FixedPointTypeClass.scala 43:59]
  wire [49:0] muls_3; // @[FixedPointTypeClass.scala 43:59]
  wire [49:0] muls_4; // @[FixedPointTypeClass.scala 43:59]
  wire [32:0] muls_5; // @[FixedPointTypeClass.scala 43:59]
  wire [48:0] _GEN_19; // @[FixedPointTypeClass.scala 21:58]
  wire [48:0] _T_8; // @[FixedPointTypeClass.scala 21:58]
  wire [48:0] accumulator_1; // @[FixedPointTypeClass.scala 21:58]
  wire [48:0] _T_10; // @[FixedPointTypeClass.scala 21:58]
  wire [48:0] accumulator_2; // @[FixedPointTypeClass.scala 21:58]
  wire [49:0] _GEN_20; // @[FixedPointTypeClass.scala 21:58]
  wire [49:0] _T_12; // @[FixedPointTypeClass.scala 21:58]
  wire [49:0] accumulator_3; // @[FixedPointTypeClass.scala 21:58]
  wire [49:0] _T_14; // @[FixedPointTypeClass.scala 21:58]
  wire [49:0] accumulator_4; // @[FixedPointTypeClass.scala 21:58]
  wire [49:0] _GEN_21; // @[FixedPointTypeClass.scala 21:58]
  wire [49:0] _T_16; // @[FixedPointTypeClass.scala 21:58]
  wire [49:0] accumulator_5; // @[FixedPointTypeClass.scala 21:58]
  reg  _T_18; // @[Reg.scala 19:20]
  reg [31:0] _RAND_6;
  reg  _T_19; // @[Reg.scala 19:20]
  reg [31:0] _RAND_7;
  reg  _T_20; // @[Reg.scala 19:20]
  reg [31:0] _RAND_8;
  reg  _T_21; // @[Reg.scala 19:20]
  reg [31:0] _RAND_9;
  reg  _T_22; // @[Reg.scala 19:20]
  reg [31:0] _RAND_10;
  reg  _T_23; // @[Reg.scala 19:20]
  reg [31:0] _RAND_11;
  wire [35:0] _GEN_22; // @[FIRFilter.scala 67:15]
  wire [31:0] _GEN_23; // @[FIRFilter.scala 67:15]
  assign accumulator_0 = $signed(regs_0) * $signed(32'sh4000); // @[FixedPointTypeClass.scala 43:59]
  assign muls_1 = $signed(regs_1) * $signed(32'sh8000); // @[FixedPointTypeClass.scala 43:59]
  assign muls_2 = $signed(regs_2) * $signed(32'shc000); // @[FixedPointTypeClass.scala 43:59]
  assign muls_3 = $signed(regs_3) * $signed(32'sh10000); // @[FixedPointTypeClass.scala 43:59]
  assign muls_4 = $signed(regs_4) * $signed(32'sh14000); // @[FixedPointTypeClass.scala 43:59]
  assign muls_5 = $signed(regs_5) * $signed(32'sh0); // @[FixedPointTypeClass.scala 43:59]
  assign _GEN_19 = {{1{accumulator_0[47]}},accumulator_0}; // @[FixedPointTypeClass.scala 21:58]
  assign _T_8 = $signed(muls_1) + $signed(_GEN_19); // @[FixedPointTypeClass.scala 21:58]
  assign accumulator_1 = $signed(_T_8); // @[FixedPointTypeClass.scala 21:58]
  assign _T_10 = $signed(muls_2) + $signed(accumulator_1); // @[FixedPointTypeClass.scala 21:58]
  assign accumulator_2 = $signed(_T_10); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_20 = {{1{accumulator_2[48]}},accumulator_2}; // @[FixedPointTypeClass.scala 21:58]
  assign _T_12 = $signed(muls_3) + $signed(_GEN_20); // @[FixedPointTypeClass.scala 21:58]
  assign accumulator_3 = $signed(_T_12); // @[FixedPointTypeClass.scala 21:58]
  assign _T_14 = $signed(muls_4) + $signed(accumulator_3); // @[FixedPointTypeClass.scala 21:58]
  assign accumulator_4 = $signed(_T_14); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_21 = {{17{muls_5[32]}},muls_5}; // @[FixedPointTypeClass.scala 21:58]
  assign _T_16 = $signed(_GEN_21) + $signed(accumulator_4); // @[FixedPointTypeClass.scala 21:58]
  assign accumulator_5 = $signed(_T_16); // @[FixedPointTypeClass.scala 21:58]
  assign io_out_valid = _T_23 & io_in_valid; // @[FIRFilter.scala 68:16]
  assign _GEN_22 = accumulator_5[49:14]; // @[FIRFilter.scala 67:15]
  assign _GEN_23 = _GEN_22[31:0]; // @[FIRFilter.scala 67:15]
  assign io_out_bits = $signed(_GEN_23); // @[FIRFilter.scala 67:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  regs_3 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  regs_4 = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  regs_5 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_18 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_19 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_20 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_21 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_22 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_23 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      regs_0 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_0 <= io_in_bits;
      end
    end
    if (reset) begin
      regs_1 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_1 <= regs_0;
      end
    end
    if (reset) begin
      regs_2 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_2 <= regs_1;
      end
    end
    if (reset) begin
      regs_3 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_3 <= regs_2;
      end
    end
    if (reset) begin
      regs_4 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_4 <= regs_3;
      end
    end
    if (reset) begin
      regs_5 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_5 <= regs_4;
      end
    end
    if (reset) begin
      _T_18 <= 1'h0;
    end else begin
      if (io_in_valid) begin
        _T_18 <= io_in_valid;
      end
    end
    if (reset) begin
      _T_19 <= 1'h0;
    end else begin
      if (io_in_valid) begin
        _T_19 <= _T_18;
      end
    end
    if (reset) begin
      _T_20 <= 1'h0;
    end else begin
      if (io_in_valid) begin
        _T_20 <= _T_19;
      end
    end
    if (reset) begin
      _T_21 <= 1'h0;
    end else begin
      if (io_in_valid) begin
        _T_21 <= _T_20;
      end
    end
    if (reset) begin
      _T_22 <= 1'h0;
    end else begin
      if (io_in_valid) begin
        _T_22 <= _T_21;
      end
    end
    if (reset) begin
      _T_23 <= 1'h0;
    end else begin
      if (io_in_valid) begin
        _T_23 <= _T_22;
      end
    end
  end
endmodule
module lineLength(
  input         clock,
  input         reset,
  input         io_in_valid,
  input  [31:0] io_in_bits,
  output        io_out_valid,
  output [31:0] io_out_bits
);
  reg [31:0] lineLengths_0; // @[lineLength.scala 47:28]
  reg [31:0] _RAND_0;
  reg [31:0] pastVal; // @[lineLength.scala 49:24]
  reg [31:0] _RAND_1;
  wire  _T_3; // @[FixedPointTypeClass.scala 57:62]
  wire [31:0] _T_5; // @[FixedPointTypeClass.scala 31:68]
  wire [31:0] _T_6; // @[FixedPointTypeClass.scala 31:68]
  wire [31:0] _T_8; // @[FixedPointTypeClass.scala 31:68]
  wire [31:0] _T_9; // @[FixedPointTypeClass.scala 31:68]
  wire [30:0] _T_12; // @[FixedPointTypeClass.scala 118:50]
  wire [27:0] _T_13; // @[FixedPointTypeClass.scala 118:50]
  reg  _T_14; // @[Reg.scala 19:20]
  reg [31:0] _RAND_2;
  reg  _T_15; // @[Reg.scala 19:20]
  reg [31:0] _RAND_3;
  assign _T_3 = $signed(io_in_bits) >= $signed(pastVal); // @[FixedPointTypeClass.scala 57:62]
  assign _T_5 = $signed(io_in_bits) - $signed(pastVal); // @[FixedPointTypeClass.scala 31:68]
  assign _T_6 = $signed(_T_5); // @[FixedPointTypeClass.scala 31:68]
  assign _T_8 = $signed(pastVal) - $signed(io_in_bits); // @[FixedPointTypeClass.scala 31:68]
  assign _T_9 = $signed(_T_8); // @[FixedPointTypeClass.scala 31:68]
  assign _T_12 = lineLengths_0[31:1]; // @[FixedPointTypeClass.scala 118:50]
  assign _T_13 = _T_12[30:3]; // @[FixedPointTypeClass.scala 118:50]
  assign io_out_valid = _T_15 & io_in_valid; // @[lineLength.scala 84:16]
  assign io_out_bits = {{4{_T_13[27]}},_T_13}; // @[lineLength.scala 83:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  lineLengths_0 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  pastVal = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_14 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_15 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      lineLengths_0 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        if (_T_3) begin
          lineLengths_0 <= _T_6;
        end else begin
          lineLengths_0 <= _T_9;
        end
      end
    end
    if (reset) begin
      pastVal <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        pastVal <= io_in_bits;
      end
    end
    if (reset) begin
      _T_14 <= 1'h0;
    end else begin
      if (io_in_valid) begin
        _T_14 <= io_in_valid;
      end
    end
    if (reset) begin
      _T_15 <= 1'h0;
    end else begin
      if (io_in_valid) begin
        _T_15 <= _T_14;
      end
    end
  end
endmodule
module sumSquares(
  input         clock,
  input         reset,
  input         io_in_valid,
  input  [31:0] io_in_bits,
  output        io_out_valid,
  output [31:0] io_out_bits
);
  reg [31:0] sumSquaress_0; // @[SumSquares.scala 41:28]
  reg [31:0] _RAND_0;
  wire [63:0] _T_3; // @[FixedPointTypeClass.scala 43:59]
  wire [39:0] _GEN_7; // @[SumSquares.scala 52:31]
  wire [39:0] _GEN_8; // @[SumSquares.scala 52:31]
  wire [63:0] _GEN_1; // @[SumSquares.scala 52:31]
  wire [30:0] _T_5; // @[FixedPointTypeClass.scala 118:50]
  wire [27:0] _T_6; // @[FixedPointTypeClass.scala 118:50]
  reg  _T_7; // @[Reg.scala 19:20]
  reg [31:0] _RAND_1;
  reg  _T_8; // @[Reg.scala 19:20]
  reg [31:0] _RAND_2;
  wire [55:0] _GEN_10; // @[SumSquares.scala 53:34 SumSquares.scala 56:22]
  wire [31:0] _GEN_11; // @[SumSquares.scala 53:34 SumSquares.scala 56:22]
  assign _T_3 = $signed(io_in_bits) * $signed(io_in_bits); // @[FixedPointTypeClass.scala 43:59]
  assign _GEN_7 = {{8{sumSquaress_0[31]}},sumSquaress_0}; // @[SumSquares.scala 52:31]
  assign _GEN_8 = $signed(_GEN_7) << 8; // @[SumSquares.scala 52:31]
  assign _GEN_1 = io_in_valid ? $signed(_T_3) : $signed({{24{_GEN_8[39]}},_GEN_8}); // @[SumSquares.scala 52:31]
  assign _T_5 = sumSquaress_0[31:1]; // @[FixedPointTypeClass.scala 118:50]
  assign _T_6 = _T_5[30:3]; // @[FixedPointTypeClass.scala 118:50]
  assign io_out_valid = _T_8 & io_in_valid; // @[SumSquares.scala 78:16]
  assign io_out_bits = {{4{_T_6[27]}},_T_6}; // @[SumSquares.scala 77:15]
  assign _GEN_10 = _GEN_1[63:8]; // @[SumSquares.scala 53:34 SumSquares.scala 56:22]
  assign _GEN_11 = _GEN_10[31:0]; // @[SumSquares.scala 53:34 SumSquares.scala 56:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sumSquaress_0 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_7 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_8 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      sumSquaress_0 <= 32'sh0;
    end else begin
      sumSquaress_0 <= $signed(_GEN_11);
    end
    if (reset) begin
      _T_7 <= 1'h0;
    end else begin
      if (io_in_valid) begin
        _T_7 <= io_in_valid;
      end
    end
    if (reset) begin
      _T_8 <= 1'h0;
    end else begin
      if (io_in_valid) begin
        _T_8 <= _T_7;
      end
    end
  end
endmodule
module NeuralNet(
  input         clock,
  input         io_in_valid,
  input  [31:0] io_in_bits_0,
  input  [31:0] io_in_bits_1,
  input  [31:0] io_in_bits_2,
  input  [31:0] io_in_bits_3,
  output        io_out_valid,
  output        io_out_bits,
  input  [31:0] io_inputWeights_0_0,
  input  [31:0] io_inputWeights_0_1,
  input  [31:0] io_inputWeights_0_2,
  input  [31:0] io_inputWeights_0_3,
  input  [31:0] io_inputWeights_1_0,
  input  [31:0] io_inputWeights_1_1,
  input  [31:0] io_inputWeights_1_2,
  input  [31:0] io_inputWeights_1_3,
  input  [31:0] io_inputWeights_2_0,
  input  [31:0] io_inputWeights_2_1,
  input  [31:0] io_inputWeights_2_2,
  input  [31:0] io_inputWeights_2_3,
  input  [31:0] io_inputWeights_3_0,
  input  [31:0] io_inputWeights_3_1,
  input  [31:0] io_inputWeights_3_2,
  input  [31:0] io_inputWeights_3_3,
  input  [31:0] io_inputWeights_4_0,
  input  [31:0] io_inputWeights_4_1,
  input  [31:0] io_inputWeights_4_2,
  input  [31:0] io_inputWeights_4_3,
  input  [31:0] io_inputWeights_5_0,
  input  [31:0] io_inputWeights_5_1,
  input  [31:0] io_inputWeights_5_2,
  input  [31:0] io_inputWeights_5_3,
  input  [31:0] io_inputWeights_6_0,
  input  [31:0] io_inputWeights_6_1,
  input  [31:0] io_inputWeights_6_2,
  input  [31:0] io_inputWeights_6_3,
  input  [31:0] io_inputWeights_7_0,
  input  [31:0] io_inputWeights_7_1,
  input  [31:0] io_inputWeights_7_2,
  input  [31:0] io_inputWeights_7_3,
  input  [31:0] io_inputWeights_8_0,
  input  [31:0] io_inputWeights_8_1,
  input  [31:0] io_inputWeights_8_2,
  input  [31:0] io_inputWeights_8_3,
  input  [31:0] io_inputWeights_9_0,
  input  [31:0] io_inputWeights_9_1,
  input  [31:0] io_inputWeights_9_2,
  input  [31:0] io_inputWeights_9_3,
  input  [31:0] io_midAndOutputWeights_0_0,
  input  [31:0] io_midAndOutputWeights_0_1,
  input  [31:0] io_midAndOutputWeights_0_2,
  input  [31:0] io_midAndOutputWeights_0_3,
  input  [31:0] io_midAndOutputWeights_0_4,
  input  [31:0] io_midAndOutputWeights_0_5,
  input  [31:0] io_midAndOutputWeights_0_6,
  input  [31:0] io_midAndOutputWeights_0_7,
  input  [31:0] io_midAndOutputWeights_0_8,
  input  [31:0] io_midAndOutputWeights_0_9,
  input  [31:0] io_midAndOutputWeights_1_0,
  input  [31:0] io_midAndOutputWeights_1_1,
  input  [31:0] io_midAndOutputWeights_1_2,
  input  [31:0] io_midAndOutputWeights_1_3,
  input  [31:0] io_midAndOutputWeights_1_4,
  input  [31:0] io_midAndOutputWeights_1_5,
  input  [31:0] io_midAndOutputWeights_1_6,
  input  [31:0] io_midAndOutputWeights_1_7,
  input  [31:0] io_midAndOutputWeights_1_8,
  input  [31:0] io_midAndOutputWeights_1_9,
  input  [31:0] io_midAndOutputWeights_2_0,
  input  [31:0] io_midAndOutputWeights_2_1,
  input  [31:0] io_midAndOutputWeights_2_2,
  input  [31:0] io_midAndOutputWeights_2_3,
  input  [31:0] io_midAndOutputWeights_2_4,
  input  [31:0] io_midAndOutputWeights_2_5,
  input  [31:0] io_midAndOutputWeights_2_6,
  input  [31:0] io_midAndOutputWeights_2_7,
  input  [31:0] io_midAndOutputWeights_2_8,
  input  [31:0] io_midAndOutputWeights_2_9,
  input  [31:0] io_midAndOutputWeights_3_0,
  input  [31:0] io_midAndOutputWeights_3_1,
  input  [31:0] io_midAndOutputWeights_3_2,
  input  [31:0] io_midAndOutputWeights_3_3,
  input  [31:0] io_midAndOutputWeights_3_4,
  input  [31:0] io_midAndOutputWeights_3_5,
  input  [31:0] io_midAndOutputWeights_3_6,
  input  [31:0] io_midAndOutputWeights_3_7,
  input  [31:0] io_midAndOutputWeights_3_8,
  input  [31:0] io_midAndOutputWeights_3_9,
  input  [31:0] io_midAndOutputWeights_4_0,
  input  [31:0] io_midAndOutputWeights_4_1,
  input  [31:0] io_midAndOutputWeights_4_2,
  input  [31:0] io_midAndOutputWeights_4_3,
  input  [31:0] io_midAndOutputWeights_4_4,
  input  [31:0] io_midAndOutputWeights_4_5,
  input  [31:0] io_midAndOutputWeights_4_6,
  input  [31:0] io_midAndOutputWeights_4_7,
  input  [31:0] io_midAndOutputWeights_4_8,
  input  [31:0] io_midAndOutputWeights_4_9,
  input  [31:0] io_midAndOutputWeights_5_0,
  input  [31:0] io_midAndOutputWeights_5_1,
  input  [31:0] io_midAndOutputWeights_5_2,
  input  [31:0] io_midAndOutputWeights_5_3,
  input  [31:0] io_midAndOutputWeights_5_4,
  input  [31:0] io_midAndOutputWeights_5_5,
  input  [31:0] io_midAndOutputWeights_5_6,
  input  [31:0] io_midAndOutputWeights_5_7,
  input  [31:0] io_midAndOutputWeights_5_8,
  input  [31:0] io_midAndOutputWeights_5_9,
  input  [31:0] io_midAndOutputWeights_6_0,
  input  [31:0] io_midAndOutputWeights_6_1,
  input  [31:0] io_midAndOutputWeights_6_2,
  input  [31:0] io_midAndOutputWeights_6_3,
  input  [31:0] io_midAndOutputWeights_6_4,
  input  [31:0] io_midAndOutputWeights_6_5,
  input  [31:0] io_midAndOutputWeights_6_6,
  input  [31:0] io_midAndOutputWeights_6_7,
  input  [31:0] io_midAndOutputWeights_6_8,
  input  [31:0] io_midAndOutputWeights_6_9,
  input  [31:0] io_midAndOutputWeights_7_0,
  input  [31:0] io_midAndOutputWeights_7_1,
  input  [31:0] io_midAndOutputWeights_7_2,
  input  [31:0] io_midAndOutputWeights_7_3,
  input  [31:0] io_midAndOutputWeights_7_4,
  input  [31:0] io_midAndOutputWeights_7_5,
  input  [31:0] io_midAndOutputWeights_7_6,
  input  [31:0] io_midAndOutputWeights_7_7,
  input  [31:0] io_midAndOutputWeights_7_8,
  input  [31:0] io_midAndOutputWeights_7_9,
  input  [31:0] io_midAndOutputWeights_8_0,
  input  [31:0] io_midAndOutputWeights_8_1,
  input  [31:0] io_midAndOutputWeights_8_2,
  input  [31:0] io_midAndOutputWeights_8_3,
  input  [31:0] io_midAndOutputWeights_8_4,
  input  [31:0] io_midAndOutputWeights_8_5,
  input  [31:0] io_midAndOutputWeights_8_6,
  input  [31:0] io_midAndOutputWeights_8_7,
  input  [31:0] io_midAndOutputWeights_8_8,
  input  [31:0] io_midAndOutputWeights_8_9,
  input  [31:0] io_midAndOutputWeights_9_0,
  input  [31:0] io_midAndOutputWeights_9_1,
  input  [31:0] io_midAndOutputWeights_9_2,
  input  [31:0] io_midAndOutputWeights_9_3,
  input  [31:0] io_midAndOutputWeights_9_4,
  input  [31:0] io_midAndOutputWeights_9_5,
  input  [31:0] io_midAndOutputWeights_9_6,
  input  [31:0] io_midAndOutputWeights_9_7,
  input  [31:0] io_midAndOutputWeights_9_8,
  input  [31:0] io_midAndOutputWeights_9_9,
  input  [31:0] io_midAndOutputWeights_10_0,
  input  [31:0] io_midAndOutputWeights_10_1,
  input  [31:0] io_midAndOutputWeights_10_2,
  input  [31:0] io_midAndOutputWeights_10_3,
  input  [31:0] io_midAndOutputWeights_10_4,
  input  [31:0] io_midAndOutputWeights_10_5,
  input  [31:0] io_midAndOutputWeights_10_6,
  input  [31:0] io_midAndOutputWeights_10_7,
  input  [31:0] io_midAndOutputWeights_10_8,
  input  [31:0] io_midAndOutputWeights_10_9,
  input  [31:0] io_midAndOutputWeights_11_0,
  input  [31:0] io_midAndOutputWeights_11_1,
  input  [31:0] io_midAndOutputWeights_11_2,
  input  [31:0] io_midAndOutputWeights_11_3,
  input  [31:0] io_midAndOutputWeights_11_4,
  input  [31:0] io_midAndOutputWeights_11_5,
  input  [31:0] io_midAndOutputWeights_11_6,
  input  [31:0] io_midAndOutputWeights_11_7,
  input  [31:0] io_midAndOutputWeights_11_8,
  input  [31:0] io_midAndOutputWeights_11_9,
  input  [31:0] io_midAndOutputWeights_12_0,
  input  [31:0] io_midAndOutputWeights_12_1,
  input  [31:0] io_midAndOutputWeights_12_2,
  input  [31:0] io_midAndOutputWeights_12_3,
  input  [31:0] io_midAndOutputWeights_12_4,
  input  [31:0] io_midAndOutputWeights_12_5,
  input  [31:0] io_midAndOutputWeights_12_6,
  input  [31:0] io_midAndOutputWeights_12_7,
  input  [31:0] io_midAndOutputWeights_12_8,
  input  [31:0] io_midAndOutputWeights_12_9,
  input  [31:0] io_midAndOutputWeights_13_0,
  input  [31:0] io_midAndOutputWeights_13_1,
  input  [31:0] io_midAndOutputWeights_13_2,
  input  [31:0] io_midAndOutputWeights_13_3,
  input  [31:0] io_midAndOutputWeights_13_4,
  input  [31:0] io_midAndOutputWeights_13_5,
  input  [31:0] io_midAndOutputWeights_13_6,
  input  [31:0] io_midAndOutputWeights_13_7,
  input  [31:0] io_midAndOutputWeights_13_8,
  input  [31:0] io_midAndOutputWeights_13_9,
  input  [31:0] io_midAndOutputWeights_14_0,
  input  [31:0] io_midAndOutputWeights_14_1,
  input  [31:0] io_midAndOutputWeights_14_2,
  input  [31:0] io_midAndOutputWeights_14_3,
  input  [31:0] io_midAndOutputWeights_14_4,
  input  [31:0] io_midAndOutputWeights_14_5,
  input  [31:0] io_midAndOutputWeights_14_6,
  input  [31:0] io_midAndOutputWeights_14_7,
  input  [31:0] io_midAndOutputWeights_14_8,
  input  [31:0] io_midAndOutputWeights_14_9,
  input  [31:0] io_midAndOutputWeights_15_0,
  input  [31:0] io_midAndOutputWeights_15_1,
  input  [31:0] io_midAndOutputWeights_15_2,
  input  [31:0] io_midAndOutputWeights_15_3,
  input  [31:0] io_midAndOutputWeights_15_4,
  input  [31:0] io_midAndOutputWeights_15_5,
  input  [31:0] io_midAndOutputWeights_15_6,
  input  [31:0] io_midAndOutputWeights_15_7,
  input  [31:0] io_midAndOutputWeights_15_8,
  input  [31:0] io_midAndOutputWeights_15_9,
  input  [31:0] io_midAndOutputWeights_16_0,
  input  [31:0] io_midAndOutputWeights_16_1,
  input  [31:0] io_midAndOutputWeights_16_2,
  input  [31:0] io_midAndOutputWeights_16_3,
  input  [31:0] io_midAndOutputWeights_16_4,
  input  [31:0] io_midAndOutputWeights_16_5,
  input  [31:0] io_midAndOutputWeights_16_6,
  input  [31:0] io_midAndOutputWeights_16_7,
  input  [31:0] io_midAndOutputWeights_16_8,
  input  [31:0] io_midAndOutputWeights_16_9,
  input  [31:0] io_midAndOutputWeights_17_0,
  input  [31:0] io_midAndOutputWeights_17_1,
  input  [31:0] io_midAndOutputWeights_17_2,
  input  [31:0] io_midAndOutputWeights_17_3,
  input  [31:0] io_midAndOutputWeights_17_4,
  input  [31:0] io_midAndOutputWeights_17_5,
  input  [31:0] io_midAndOutputWeights_17_6,
  input  [31:0] io_midAndOutputWeights_17_7,
  input  [31:0] io_midAndOutputWeights_17_8,
  input  [31:0] io_midAndOutputWeights_17_9,
  input  [31:0] io_midAndOutputWeights_18_0,
  input  [31:0] io_midAndOutputWeights_18_1,
  input  [31:0] io_midAndOutputWeights_18_2,
  input  [31:0] io_midAndOutputWeights_18_3,
  input  [31:0] io_midAndOutputWeights_18_4,
  input  [31:0] io_midAndOutputWeights_18_5,
  input  [31:0] io_midAndOutputWeights_18_6,
  input  [31:0] io_midAndOutputWeights_18_7,
  input  [31:0] io_midAndOutputWeights_18_8,
  input  [31:0] io_midAndOutputWeights_18_9,
  input  [31:0] io_midAndOutputWeights_19_0,
  input  [31:0] io_midAndOutputWeights_19_1,
  input  [31:0] io_midAndOutputWeights_19_2,
  input  [31:0] io_midAndOutputWeights_19_3,
  input  [31:0] io_midAndOutputWeights_19_4,
  input  [31:0] io_midAndOutputWeights_19_5,
  input  [31:0] io_midAndOutputWeights_19_6,
  input  [31:0] io_midAndOutputWeights_19_7,
  input  [31:0] io_midAndOutputWeights_19_8,
  input  [31:0] io_midAndOutputWeights_19_9,
  input  [31:0] io_midAndOutputWeights_20_0,
  input  [31:0] io_midAndOutputWeights_20_1,
  input  [31:0] io_midAndOutputWeights_20_2,
  input  [31:0] io_midAndOutputWeights_20_3,
  input  [31:0] io_midAndOutputWeights_20_4,
  input  [31:0] io_midAndOutputWeights_20_5,
  input  [31:0] io_midAndOutputWeights_20_6,
  input  [31:0] io_midAndOutputWeights_20_7,
  input  [31:0] io_midAndOutputWeights_20_8,
  input  [31:0] io_midAndOutputWeights_20_9,
  input  [31:0] io_biasVecs_0_0,
  input  [31:0] io_biasVecs_0_1,
  input  [31:0] io_biasVecs_0_2,
  input  [31:0] io_biasVecs_0_3,
  input  [31:0] io_biasVecs_0_4,
  input  [31:0] io_biasVecs_0_5,
  input  [31:0] io_biasVecs_0_6,
  input  [31:0] io_biasVecs_0_7,
  input  [31:0] io_biasVecs_0_8,
  input  [31:0] io_biasVecs_0_9,
  input  [31:0] io_biasVecs_1_0,
  input  [31:0] io_biasVecs_1_1,
  input  [31:0] io_biasVecs_1_2,
  input  [31:0] io_biasVecs_1_3,
  input  [31:0] io_biasVecs_1_4,
  input  [31:0] io_biasVecs_1_5,
  input  [31:0] io_biasVecs_1_6,
  input  [31:0] io_biasVecs_1_7,
  input  [31:0] io_biasVecs_1_8,
  input  [31:0] io_biasVecs_1_9,
  input  [31:0] io_biasVecs_2_0,
  input  [31:0] io_biasVecs_2_1,
  input  [31:0] io_biasVecs_2_2,
  input  [31:0] io_biasVecs_2_3,
  input  [31:0] io_biasVecs_2_4,
  input  [31:0] io_biasVecs_2_5,
  input  [31:0] io_biasVecs_2_6,
  input  [31:0] io_biasVecs_2_7,
  input  [31:0] io_biasVecs_2_8,
  input  [31:0] io_biasVecs_2_9,
  input  [31:0] io_outputBias,
  output [31:0] io_rawVotes
);
  wire [63:0] _T; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_2; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_3; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_5; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_6; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_8; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_9; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_11; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_12; // @[FixedPointTypeClass.scala 21:58]
  wire [39:0] _GEN_2; // @[FixedPointTypeClass.scala 21:58]
  wire [39:0] _GEN_3; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _GEN_4; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_14; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_15; // @[FixedPointTypeClass.scala 21:58]
  wire  _T_16; // @[FixedPointTypeClass.scala 56:59]
  wire [63:0] _T_17; // @[neuralNet.scala 50:30]
  wire [63:0] _T_18; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_19; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_20; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_21; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_23; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_24; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_26; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_27; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_29; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_30; // @[FixedPointTypeClass.scala 21:58]
  wire [39:0] _GEN_5; // @[FixedPointTypeClass.scala 21:58]
  wire [39:0] _GEN_6; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _GEN_7; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_32; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_33; // @[FixedPointTypeClass.scala 21:58]
  wire  _T_34; // @[FixedPointTypeClass.scala 56:59]
  wire [63:0] _T_35; // @[neuralNet.scala 50:30]
  wire [63:0] _T_36; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_37; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_38; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_39; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_41; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_42; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_44; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_45; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_47; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_48; // @[FixedPointTypeClass.scala 21:58]
  wire [39:0] _GEN_8; // @[FixedPointTypeClass.scala 21:58]
  wire [39:0] _GEN_9; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _GEN_10; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_50; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_51; // @[FixedPointTypeClass.scala 21:58]
  wire  _T_52; // @[FixedPointTypeClass.scala 56:59]
  wire [63:0] _T_53; // @[neuralNet.scala 50:30]
  wire [63:0] _T_54; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_55; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_56; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_57; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_59; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_60; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_62; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_63; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_65; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_66; // @[FixedPointTypeClass.scala 21:58]
  wire [39:0] _GEN_11; // @[FixedPointTypeClass.scala 21:58]
  wire [39:0] _GEN_12; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _GEN_13; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_68; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_69; // @[FixedPointTypeClass.scala 21:58]
  wire  _T_70; // @[FixedPointTypeClass.scala 56:59]
  wire [63:0] _T_71; // @[neuralNet.scala 50:30]
  wire [63:0] _T_72; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_73; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_74; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_75; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_77; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_78; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_80; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_81; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_83; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_84; // @[FixedPointTypeClass.scala 21:58]
  wire [39:0] _GEN_14; // @[FixedPointTypeClass.scala 21:58]
  wire [39:0] _GEN_15; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _GEN_16; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_86; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_87; // @[FixedPointTypeClass.scala 21:58]
  wire  _T_88; // @[FixedPointTypeClass.scala 56:59]
  wire [63:0] _T_89; // @[neuralNet.scala 50:30]
  wire [63:0] _T_90; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_91; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_92; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_93; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_95; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_96; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_98; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_99; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_101; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_102; // @[FixedPointTypeClass.scala 21:58]
  wire [39:0] _GEN_17; // @[FixedPointTypeClass.scala 21:58]
  wire [39:0] _GEN_18; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _GEN_19; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_104; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_105; // @[FixedPointTypeClass.scala 21:58]
  wire  _T_106; // @[FixedPointTypeClass.scala 56:59]
  wire [63:0] _T_107; // @[neuralNet.scala 50:30]
  wire [63:0] _T_108; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_109; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_110; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_111; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_113; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_114; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_116; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_117; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_119; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_120; // @[FixedPointTypeClass.scala 21:58]
  wire [39:0] _GEN_20; // @[FixedPointTypeClass.scala 21:58]
  wire [39:0] _GEN_21; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _GEN_22; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_122; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_123; // @[FixedPointTypeClass.scala 21:58]
  wire  _T_124; // @[FixedPointTypeClass.scala 56:59]
  wire [63:0] _T_125; // @[neuralNet.scala 50:30]
  wire [63:0] _T_126; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_127; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_128; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_129; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_131; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_132; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_134; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_135; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_137; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_138; // @[FixedPointTypeClass.scala 21:58]
  wire [39:0] _GEN_23; // @[FixedPointTypeClass.scala 21:58]
  wire [39:0] _GEN_24; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _GEN_25; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_140; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_141; // @[FixedPointTypeClass.scala 21:58]
  wire  _T_142; // @[FixedPointTypeClass.scala 56:59]
  wire [63:0] _T_143; // @[neuralNet.scala 50:30]
  wire [63:0] _T_144; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_145; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_146; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_147; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_149; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_150; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_152; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_153; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_155; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_156; // @[FixedPointTypeClass.scala 21:58]
  wire [39:0] _GEN_26; // @[FixedPointTypeClass.scala 21:58]
  wire [39:0] _GEN_27; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _GEN_28; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_158; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_159; // @[FixedPointTypeClass.scala 21:58]
  wire  _T_160; // @[FixedPointTypeClass.scala 56:59]
  wire [63:0] _T_161; // @[neuralNet.scala 50:30]
  wire [63:0] _T_162; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_163; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_164; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_165; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_167; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_168; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_170; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_171; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_173; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_174; // @[FixedPointTypeClass.scala 21:58]
  wire [39:0] _GEN_29; // @[FixedPointTypeClass.scala 21:58]
  wire [39:0] _GEN_30; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _GEN_31; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_176; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_177; // @[FixedPointTypeClass.scala 21:58]
  wire  _T_178; // @[FixedPointTypeClass.scala 56:59]
  wire [63:0] _T_179; // @[neuralNet.scala 50:30]
  wire [55:0] _GEN_32; // @[neuralNet.scala 43:26 neuralNet.scala 50:24]
  wire [31:0] _GEN_33; // @[neuralNet.scala 43:26 neuralNet.scala 50:24]
  wire [31:0] hiddenLayers_0_0; // @[neuralNet.scala 43:26 neuralNet.scala 50:24]
  wire [63:0] _T_180; // @[FixedPointTypeClass.scala 43:59]
  wire [55:0] _GEN_34; // @[neuralNet.scala 43:26 neuralNet.scala 50:24]
  wire [31:0] _GEN_35; // @[neuralNet.scala 43:26 neuralNet.scala 50:24]
  wire [31:0] hiddenLayers_0_1; // @[neuralNet.scala 43:26 neuralNet.scala 50:24]
  wire [63:0] _T_181; // @[FixedPointTypeClass.scala 43:59]
  wire [55:0] _GEN_36; // @[neuralNet.scala 43:26 neuralNet.scala 50:24]
  wire [31:0] _GEN_37; // @[neuralNet.scala 43:26 neuralNet.scala 50:24]
  wire [31:0] hiddenLayers_0_2; // @[neuralNet.scala 43:26 neuralNet.scala 50:24]
  wire [63:0] _T_182; // @[FixedPointTypeClass.scala 43:59]
  wire [55:0] _GEN_38; // @[neuralNet.scala 43:26 neuralNet.scala 50:24]
  wire [31:0] _GEN_39; // @[neuralNet.scala 43:26 neuralNet.scala 50:24]
  wire [31:0] hiddenLayers_0_3; // @[neuralNet.scala 43:26 neuralNet.scala 50:24]
  wire [63:0] _T_183; // @[FixedPointTypeClass.scala 43:59]
  wire [55:0] _GEN_40; // @[neuralNet.scala 43:26 neuralNet.scala 50:24]
  wire [31:0] _GEN_41; // @[neuralNet.scala 43:26 neuralNet.scala 50:24]
  wire [31:0] hiddenLayers_0_4; // @[neuralNet.scala 43:26 neuralNet.scala 50:24]
  wire [63:0] _T_184; // @[FixedPointTypeClass.scala 43:59]
  wire [55:0] _GEN_42; // @[neuralNet.scala 43:26 neuralNet.scala 50:24]
  wire [31:0] _GEN_43; // @[neuralNet.scala 43:26 neuralNet.scala 50:24]
  wire [31:0] hiddenLayers_0_5; // @[neuralNet.scala 43:26 neuralNet.scala 50:24]
  wire [63:0] _T_185; // @[FixedPointTypeClass.scala 43:59]
  wire [55:0] _GEN_44; // @[neuralNet.scala 43:26 neuralNet.scala 50:24]
  wire [31:0] _GEN_45; // @[neuralNet.scala 43:26 neuralNet.scala 50:24]
  wire [31:0] hiddenLayers_0_6; // @[neuralNet.scala 43:26 neuralNet.scala 50:24]
  wire [63:0] _T_186; // @[FixedPointTypeClass.scala 43:59]
  wire [55:0] _GEN_46; // @[neuralNet.scala 43:26 neuralNet.scala 50:24]
  wire [31:0] _GEN_47; // @[neuralNet.scala 43:26 neuralNet.scala 50:24]
  wire [31:0] hiddenLayers_0_7; // @[neuralNet.scala 43:26 neuralNet.scala 50:24]
  wire [63:0] _T_187; // @[FixedPointTypeClass.scala 43:59]
  wire [55:0] _GEN_48; // @[neuralNet.scala 43:26 neuralNet.scala 50:24]
  wire [31:0] _GEN_49; // @[neuralNet.scala 43:26 neuralNet.scala 50:24]
  wire [31:0] hiddenLayers_0_8; // @[neuralNet.scala 43:26 neuralNet.scala 50:24]
  wire [63:0] _T_188; // @[FixedPointTypeClass.scala 43:59]
  wire [55:0] _GEN_50; // @[neuralNet.scala 43:26 neuralNet.scala 50:24]
  wire [31:0] _GEN_51; // @[neuralNet.scala 43:26 neuralNet.scala 50:24]
  wire [31:0] hiddenLayers_0_9; // @[neuralNet.scala 43:26 neuralNet.scala 50:24]
  wire [63:0] _T_189; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_191; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_192; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_194; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_195; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_197; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_198; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_200; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_201; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_203; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_204; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_206; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_207; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_209; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_210; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_212; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_213; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_215; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_216; // @[FixedPointTypeClass.scala 21:58]
  wire [39:0] _GEN_52; // @[FixedPointTypeClass.scala 21:58]
  wire [39:0] _GEN_53; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _GEN_54; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_218; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_219; // @[FixedPointTypeClass.scala 21:58]
  wire  _T_220; // @[FixedPointTypeClass.scala 56:59]
  wire [63:0] _T_221; // @[neuralNet.scala 59:32]
  wire [63:0] _T_222; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_223; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_224; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_225; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_226; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_227; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_228; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_229; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_230; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_231; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_233; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_234; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_236; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_237; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_239; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_240; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_242; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_243; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_245; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_246; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_248; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_249; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_251; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_252; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_254; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_255; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_257; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_258; // @[FixedPointTypeClass.scala 21:58]
  wire [39:0] _GEN_55; // @[FixedPointTypeClass.scala 21:58]
  wire [39:0] _GEN_56; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _GEN_57; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_260; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_261; // @[FixedPointTypeClass.scala 21:58]
  wire  _T_262; // @[FixedPointTypeClass.scala 56:59]
  wire [63:0] _T_263; // @[neuralNet.scala 59:32]
  wire [63:0] _T_264; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_265; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_266; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_267; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_268; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_269; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_270; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_271; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_272; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_273; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_275; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_276; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_278; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_279; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_281; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_282; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_284; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_285; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_287; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_288; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_290; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_291; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_293; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_294; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_296; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_297; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_299; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_300; // @[FixedPointTypeClass.scala 21:58]
  wire [39:0] _GEN_58; // @[FixedPointTypeClass.scala 21:58]
  wire [39:0] _GEN_59; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _GEN_60; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_302; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_303; // @[FixedPointTypeClass.scala 21:58]
  wire  _T_304; // @[FixedPointTypeClass.scala 56:59]
  wire [63:0] _T_305; // @[neuralNet.scala 59:32]
  wire [63:0] _T_306; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_307; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_308; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_309; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_310; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_311; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_312; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_313; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_314; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_315; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_317; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_318; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_320; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_321; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_323; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_324; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_326; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_327; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_329; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_330; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_332; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_333; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_335; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_336; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_338; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_339; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_341; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_342; // @[FixedPointTypeClass.scala 21:58]
  wire [39:0] _GEN_61; // @[FixedPointTypeClass.scala 21:58]
  wire [39:0] _GEN_62; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _GEN_63; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_344; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_345; // @[FixedPointTypeClass.scala 21:58]
  wire  _T_346; // @[FixedPointTypeClass.scala 56:59]
  wire [63:0] _T_347; // @[neuralNet.scala 59:32]
  wire [63:0] _T_348; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_349; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_350; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_351; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_352; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_353; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_354; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_355; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_356; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_357; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_359; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_360; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_362; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_363; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_365; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_366; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_368; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_369; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_371; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_372; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_374; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_375; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_377; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_378; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_380; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_381; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_383; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_384; // @[FixedPointTypeClass.scala 21:58]
  wire [39:0] _GEN_64; // @[FixedPointTypeClass.scala 21:58]
  wire [39:0] _GEN_65; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _GEN_66; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_386; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_387; // @[FixedPointTypeClass.scala 21:58]
  wire  _T_388; // @[FixedPointTypeClass.scala 56:59]
  wire [63:0] _T_389; // @[neuralNet.scala 59:32]
  wire [63:0] _T_390; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_391; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_392; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_393; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_394; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_395; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_396; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_397; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_398; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_399; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_401; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_402; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_404; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_405; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_407; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_408; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_410; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_411; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_413; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_414; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_416; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_417; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_419; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_420; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_422; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_423; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_425; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_426; // @[FixedPointTypeClass.scala 21:58]
  wire [39:0] _GEN_67; // @[FixedPointTypeClass.scala 21:58]
  wire [39:0] _GEN_68; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _GEN_69; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_428; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_429; // @[FixedPointTypeClass.scala 21:58]
  wire  _T_430; // @[FixedPointTypeClass.scala 56:59]
  wire [63:0] _T_431; // @[neuralNet.scala 59:32]
  wire [63:0] _T_432; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_433; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_434; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_435; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_436; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_437; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_438; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_439; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_440; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_441; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_443; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_444; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_446; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_447; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_449; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_450; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_452; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_453; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_455; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_456; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_458; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_459; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_461; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_462; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_464; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_465; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_467; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_468; // @[FixedPointTypeClass.scala 21:58]
  wire [39:0] _GEN_70; // @[FixedPointTypeClass.scala 21:58]
  wire [39:0] _GEN_71; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _GEN_72; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_470; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_471; // @[FixedPointTypeClass.scala 21:58]
  wire  _T_472; // @[FixedPointTypeClass.scala 56:59]
  wire [63:0] _T_473; // @[neuralNet.scala 59:32]
  wire [63:0] _T_474; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_475; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_476; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_477; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_478; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_479; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_480; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_481; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_482; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_483; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_485; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_486; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_488; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_489; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_491; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_492; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_494; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_495; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_497; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_498; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_500; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_501; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_503; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_504; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_506; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_507; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_509; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_510; // @[FixedPointTypeClass.scala 21:58]
  wire [39:0] _GEN_73; // @[FixedPointTypeClass.scala 21:58]
  wire [39:0] _GEN_74; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _GEN_75; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_512; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_513; // @[FixedPointTypeClass.scala 21:58]
  wire  _T_514; // @[FixedPointTypeClass.scala 56:59]
  wire [63:0] _T_515; // @[neuralNet.scala 59:32]
  wire [63:0] _T_516; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_517; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_518; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_519; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_520; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_521; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_522; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_523; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_524; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_525; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_527; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_528; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_530; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_531; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_533; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_534; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_536; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_537; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_539; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_540; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_542; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_543; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_545; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_546; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_548; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_549; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_551; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_552; // @[FixedPointTypeClass.scala 21:58]
  wire [39:0] _GEN_76; // @[FixedPointTypeClass.scala 21:58]
  wire [39:0] _GEN_77; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _GEN_78; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_554; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_555; // @[FixedPointTypeClass.scala 21:58]
  wire  _T_556; // @[FixedPointTypeClass.scala 56:59]
  wire [63:0] _T_557; // @[neuralNet.scala 59:32]
  wire [63:0] _T_558; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_559; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_560; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_561; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_562; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_563; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_564; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_565; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_566; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_567; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_569; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_570; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_572; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_573; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_575; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_576; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_578; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_579; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_581; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_582; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_584; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_585; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_587; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_588; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_590; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_591; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_593; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_594; // @[FixedPointTypeClass.scala 21:58]
  wire [39:0] _GEN_79; // @[FixedPointTypeClass.scala 21:58]
  wire [39:0] _GEN_80; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _GEN_81; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_596; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_597; // @[FixedPointTypeClass.scala 21:58]
  wire  _T_598; // @[FixedPointTypeClass.scala 56:59]
  wire [63:0] _T_599; // @[neuralNet.scala 59:32]
  wire [55:0] _GEN_82; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  wire [31:0] _GEN_83; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  wire [31:0] hiddenLayers_1_0; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  wire [63:0] _T_600; // @[FixedPointTypeClass.scala 43:59]
  wire [55:0] _GEN_84; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  wire [31:0] _GEN_85; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  wire [31:0] hiddenLayers_1_1; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  wire [63:0] _T_601; // @[FixedPointTypeClass.scala 43:59]
  wire [55:0] _GEN_86; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  wire [31:0] _GEN_87; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  wire [31:0] hiddenLayers_1_2; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  wire [63:0] _T_602; // @[FixedPointTypeClass.scala 43:59]
  wire [55:0] _GEN_88; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  wire [31:0] _GEN_89; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  wire [31:0] hiddenLayers_1_3; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  wire [63:0] _T_603; // @[FixedPointTypeClass.scala 43:59]
  wire [55:0] _GEN_90; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  wire [31:0] _GEN_91; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  wire [31:0] hiddenLayers_1_4; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  wire [63:0] _T_604; // @[FixedPointTypeClass.scala 43:59]
  wire [55:0] _GEN_92; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  wire [31:0] _GEN_93; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  wire [31:0] hiddenLayers_1_5; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  wire [63:0] _T_605; // @[FixedPointTypeClass.scala 43:59]
  wire [55:0] _GEN_94; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  wire [31:0] _GEN_95; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  wire [31:0] hiddenLayers_1_6; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  wire [63:0] _T_606; // @[FixedPointTypeClass.scala 43:59]
  wire [55:0] _GEN_96; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  wire [31:0] _GEN_97; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  wire [31:0] hiddenLayers_1_7; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  wire [63:0] _T_607; // @[FixedPointTypeClass.scala 43:59]
  wire [55:0] _GEN_98; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  wire [31:0] _GEN_99; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  wire [31:0] hiddenLayers_1_8; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  wire [63:0] _T_608; // @[FixedPointTypeClass.scala 43:59]
  wire [55:0] _GEN_100; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  wire [31:0] _GEN_101; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  wire [31:0] hiddenLayers_1_9; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  wire [63:0] _T_609; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_611; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_612; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_614; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_615; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_617; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_618; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_620; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_621; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_623; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_624; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_626; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_627; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_629; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_630; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_632; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_633; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_635; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_636; // @[FixedPointTypeClass.scala 21:58]
  wire [39:0] _GEN_102; // @[FixedPointTypeClass.scala 21:58]
  wire [39:0] _GEN_103; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _GEN_104; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_638; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_639; // @[FixedPointTypeClass.scala 21:58]
  wire  _T_640; // @[FixedPointTypeClass.scala 56:59]
  wire [63:0] _T_641; // @[neuralNet.scala 59:32]
  wire [63:0] _T_642; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_643; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_644; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_645; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_646; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_647; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_648; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_649; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_650; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_651; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_653; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_654; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_656; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_657; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_659; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_660; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_662; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_663; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_665; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_666; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_668; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_669; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_671; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_672; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_674; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_675; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_677; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_678; // @[FixedPointTypeClass.scala 21:58]
  wire [39:0] _GEN_105; // @[FixedPointTypeClass.scala 21:58]
  wire [39:0] _GEN_106; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _GEN_107; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_680; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_681; // @[FixedPointTypeClass.scala 21:58]
  wire  _T_682; // @[FixedPointTypeClass.scala 56:59]
  wire [63:0] _T_683; // @[neuralNet.scala 59:32]
  wire [63:0] _T_684; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_685; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_686; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_687; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_688; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_689; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_690; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_691; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_692; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_693; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_695; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_696; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_698; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_699; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_701; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_702; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_704; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_705; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_707; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_708; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_710; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_711; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_713; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_714; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_716; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_717; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_719; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_720; // @[FixedPointTypeClass.scala 21:58]
  wire [39:0] _GEN_108; // @[FixedPointTypeClass.scala 21:58]
  wire [39:0] _GEN_109; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _GEN_110; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_722; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_723; // @[FixedPointTypeClass.scala 21:58]
  wire  _T_724; // @[FixedPointTypeClass.scala 56:59]
  wire [63:0] _T_725; // @[neuralNet.scala 59:32]
  wire [63:0] _T_726; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_727; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_728; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_729; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_730; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_731; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_732; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_733; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_734; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_735; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_737; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_738; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_740; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_741; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_743; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_744; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_746; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_747; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_749; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_750; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_752; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_753; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_755; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_756; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_758; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_759; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_761; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_762; // @[FixedPointTypeClass.scala 21:58]
  wire [39:0] _GEN_111; // @[FixedPointTypeClass.scala 21:58]
  wire [39:0] _GEN_112; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _GEN_113; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_764; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_765; // @[FixedPointTypeClass.scala 21:58]
  wire  _T_766; // @[FixedPointTypeClass.scala 56:59]
  wire [63:0] _T_767; // @[neuralNet.scala 59:32]
  wire [63:0] _T_768; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_769; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_770; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_771; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_772; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_773; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_774; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_775; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_776; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_777; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_779; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_780; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_782; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_783; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_785; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_786; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_788; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_789; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_791; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_792; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_794; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_795; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_797; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_798; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_800; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_801; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_803; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_804; // @[FixedPointTypeClass.scala 21:58]
  wire [39:0] _GEN_114; // @[FixedPointTypeClass.scala 21:58]
  wire [39:0] _GEN_115; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _GEN_116; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_806; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_807; // @[FixedPointTypeClass.scala 21:58]
  wire  _T_808; // @[FixedPointTypeClass.scala 56:59]
  wire [63:0] _T_809; // @[neuralNet.scala 59:32]
  wire [63:0] _T_810; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_811; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_812; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_813; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_814; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_815; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_816; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_817; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_818; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_819; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_821; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_822; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_824; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_825; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_827; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_828; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_830; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_831; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_833; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_834; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_836; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_837; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_839; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_840; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_842; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_843; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_845; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_846; // @[FixedPointTypeClass.scala 21:58]
  wire [39:0] _GEN_117; // @[FixedPointTypeClass.scala 21:58]
  wire [39:0] _GEN_118; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _GEN_119; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_848; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_849; // @[FixedPointTypeClass.scala 21:58]
  wire  _T_850; // @[FixedPointTypeClass.scala 56:59]
  wire [63:0] _T_851; // @[neuralNet.scala 59:32]
  wire [63:0] _T_852; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_853; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_854; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_855; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_856; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_857; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_858; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_859; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_860; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_861; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_863; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_864; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_866; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_867; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_869; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_870; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_872; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_873; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_875; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_876; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_878; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_879; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_881; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_882; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_884; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_885; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_887; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_888; // @[FixedPointTypeClass.scala 21:58]
  wire [39:0] _GEN_120; // @[FixedPointTypeClass.scala 21:58]
  wire [39:0] _GEN_121; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _GEN_122; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_890; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_891; // @[FixedPointTypeClass.scala 21:58]
  wire  _T_892; // @[FixedPointTypeClass.scala 56:59]
  wire [63:0] _T_893; // @[neuralNet.scala 59:32]
  wire [63:0] _T_894; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_895; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_896; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_897; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_898; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_899; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_900; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_901; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_902; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_903; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_905; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_906; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_908; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_909; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_911; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_912; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_914; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_915; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_917; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_918; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_920; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_921; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_923; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_924; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_926; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_927; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_929; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_930; // @[FixedPointTypeClass.scala 21:58]
  wire [39:0] _GEN_123; // @[FixedPointTypeClass.scala 21:58]
  wire [39:0] _GEN_124; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _GEN_125; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_932; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_933; // @[FixedPointTypeClass.scala 21:58]
  wire  _T_934; // @[FixedPointTypeClass.scala 56:59]
  wire [63:0] _T_935; // @[neuralNet.scala 59:32]
  wire [63:0] _T_936; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_937; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_938; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_939; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_940; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_941; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_942; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_943; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_944; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_945; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_947; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_948; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_950; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_951; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_953; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_954; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_956; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_957; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_959; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_960; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_962; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_963; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_965; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_966; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_968; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_969; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_971; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_972; // @[FixedPointTypeClass.scala 21:58]
  wire [39:0] _GEN_126; // @[FixedPointTypeClass.scala 21:58]
  wire [39:0] _GEN_127; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _GEN_128; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_974; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_975; // @[FixedPointTypeClass.scala 21:58]
  wire  _T_976; // @[FixedPointTypeClass.scala 56:59]
  wire [63:0] _T_977; // @[neuralNet.scala 59:32]
  wire [63:0] _T_978; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_979; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_980; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_981; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_982; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_983; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_984; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_985; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_986; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_987; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_989; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_990; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_992; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_993; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_995; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_996; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_998; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_999; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1001; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1002; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1004; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1005; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1007; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1008; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1010; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1011; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1013; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1014; // @[FixedPointTypeClass.scala 21:58]
  wire [39:0] _GEN_129; // @[FixedPointTypeClass.scala 21:58]
  wire [39:0] _GEN_130; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _GEN_131; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1016; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1017; // @[FixedPointTypeClass.scala 21:58]
  wire  _T_1018; // @[FixedPointTypeClass.scala 56:59]
  wire [63:0] _T_1019; // @[neuralNet.scala 59:32]
  wire [55:0] _GEN_132; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  wire [31:0] _GEN_133; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  wire [31:0] hiddenLayers_2_0; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  wire [63:0] _T_1020; // @[FixedPointTypeClass.scala 43:59]
  wire [55:0] _GEN_134; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  wire [31:0] _GEN_135; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  wire [31:0] hiddenLayers_2_1; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  wire [63:0] _T_1021; // @[FixedPointTypeClass.scala 43:59]
  wire [55:0] _GEN_136; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  wire [31:0] _GEN_137; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  wire [31:0] hiddenLayers_2_2; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  wire [63:0] _T_1022; // @[FixedPointTypeClass.scala 43:59]
  wire [55:0] _GEN_138; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  wire [31:0] _GEN_139; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  wire [31:0] hiddenLayers_2_3; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  wire [63:0] _T_1023; // @[FixedPointTypeClass.scala 43:59]
  wire [55:0] _GEN_140; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  wire [31:0] _GEN_141; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  wire [31:0] hiddenLayers_2_4; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  wire [63:0] _T_1024; // @[FixedPointTypeClass.scala 43:59]
  wire [55:0] _GEN_142; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  wire [31:0] _GEN_143; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  wire [31:0] hiddenLayers_2_5; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  wire [63:0] _T_1025; // @[FixedPointTypeClass.scala 43:59]
  wire [55:0] _GEN_144; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  wire [31:0] _GEN_145; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  wire [31:0] hiddenLayers_2_6; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  wire [63:0] _T_1026; // @[FixedPointTypeClass.scala 43:59]
  wire [55:0] _GEN_146; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  wire [31:0] _GEN_147; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  wire [31:0] hiddenLayers_2_7; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  wire [63:0] _T_1027; // @[FixedPointTypeClass.scala 43:59]
  wire [55:0] _GEN_148; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  wire [31:0] _GEN_149; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  wire [31:0] hiddenLayers_2_8; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  wire [63:0] _T_1028; // @[FixedPointTypeClass.scala 43:59]
  wire [55:0] _GEN_150; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  wire [31:0] _GEN_151; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  wire [31:0] hiddenLayers_2_9; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  wire [63:0] _T_1029; // @[FixedPointTypeClass.scala 43:59]
  wire [63:0] _T_1031; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1032; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1034; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1035; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1037; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1038; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1040; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1041; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1043; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1044; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1046; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1047; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1049; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1050; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1052; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1053; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1055; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1056; // @[FixedPointTypeClass.scala 21:58]
  wire [39:0] _GEN_152; // @[FixedPointTypeClass.scala 21:58]
  wire [39:0] _GEN_153; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _GEN_154; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] _T_1058; // @[FixedPointTypeClass.scala 21:58]
  wire [63:0] linearOut; // @[FixedPointTypeClass.scala 21:58]
  wire  _T_1059; // @[FixedPointTypeClass.scala 56:59]
  wire [63:0] actualVotes; // @[neuralNet.scala 69:24]
  wire  finalPredict; // @[FixedPointTypeClass.scala 56:59]
  reg [63:0] rawVotesReg; // @[Reg.scala 11:16]
  reg [63:0] _RAND_0;
  reg  outReg; // @[Reg.scala 11:16]
  reg [31:0] _RAND_1;
  reg  valReg; // @[neuralNet.scala 75:23]
  reg [31:0] _RAND_2;
  wire [55:0] _GEN_155; // @[neuralNet.scala 79:15]
  wire [31:0] _GEN_156; // @[neuralNet.scala 79:15]
  assign _T = $signed(io_in_bits_0) * $signed(io_inputWeights_0_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1 = $signed(io_in_bits_1) * $signed(io_inputWeights_0_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_2 = $signed(io_in_bits_2) * $signed(io_inputWeights_0_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_3 = $signed(io_in_bits_3) * $signed(io_inputWeights_0_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_5 = $signed(_T) + $signed(_T_1); // @[FixedPointTypeClass.scala 21:58]
  assign _T_6 = $signed(_T_5); // @[FixedPointTypeClass.scala 21:58]
  assign _T_8 = $signed(_T_6) + $signed(_T_2); // @[FixedPointTypeClass.scala 21:58]
  assign _T_9 = $signed(_T_8); // @[FixedPointTypeClass.scala 21:58]
  assign _T_11 = $signed(_T_9) + $signed(_T_3); // @[FixedPointTypeClass.scala 21:58]
  assign _T_12 = $signed(_T_11); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_2 = {{8{io_biasVecs_0_0[31]}},io_biasVecs_0_0}; // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_3 = $signed(_GEN_2) << 8; // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_4 = {{24{_GEN_3[39]}},_GEN_3}; // @[FixedPointTypeClass.scala 21:58]
  assign _T_14 = $signed(_T_12) + $signed(_GEN_4); // @[FixedPointTypeClass.scala 21:58]
  assign _T_15 = $signed(_T_14); // @[FixedPointTypeClass.scala 21:58]
  assign _T_16 = $signed(_T_15) > $signed(64'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign _T_17 = _T_16 ? $signed(_T_15) : $signed(64'sh0); // @[neuralNet.scala 50:30]
  assign _T_18 = $signed(io_in_bits_0) * $signed(io_inputWeights_1_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_19 = $signed(io_in_bits_1) * $signed(io_inputWeights_1_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_20 = $signed(io_in_bits_2) * $signed(io_inputWeights_1_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_21 = $signed(io_in_bits_3) * $signed(io_inputWeights_1_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_23 = $signed(_T_18) + $signed(_T_19); // @[FixedPointTypeClass.scala 21:58]
  assign _T_24 = $signed(_T_23); // @[FixedPointTypeClass.scala 21:58]
  assign _T_26 = $signed(_T_24) + $signed(_T_20); // @[FixedPointTypeClass.scala 21:58]
  assign _T_27 = $signed(_T_26); // @[FixedPointTypeClass.scala 21:58]
  assign _T_29 = $signed(_T_27) + $signed(_T_21); // @[FixedPointTypeClass.scala 21:58]
  assign _T_30 = $signed(_T_29); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_5 = {{8{io_biasVecs_0_1[31]}},io_biasVecs_0_1}; // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_6 = $signed(_GEN_5) << 8; // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_7 = {{24{_GEN_6[39]}},_GEN_6}; // @[FixedPointTypeClass.scala 21:58]
  assign _T_32 = $signed(_T_30) + $signed(_GEN_7); // @[FixedPointTypeClass.scala 21:58]
  assign _T_33 = $signed(_T_32); // @[FixedPointTypeClass.scala 21:58]
  assign _T_34 = $signed(_T_33) > $signed(64'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign _T_35 = _T_34 ? $signed(_T_33) : $signed(64'sh0); // @[neuralNet.scala 50:30]
  assign _T_36 = $signed(io_in_bits_0) * $signed(io_inputWeights_2_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_37 = $signed(io_in_bits_1) * $signed(io_inputWeights_2_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_38 = $signed(io_in_bits_2) * $signed(io_inputWeights_2_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_39 = $signed(io_in_bits_3) * $signed(io_inputWeights_2_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_41 = $signed(_T_36) + $signed(_T_37); // @[FixedPointTypeClass.scala 21:58]
  assign _T_42 = $signed(_T_41); // @[FixedPointTypeClass.scala 21:58]
  assign _T_44 = $signed(_T_42) + $signed(_T_38); // @[FixedPointTypeClass.scala 21:58]
  assign _T_45 = $signed(_T_44); // @[FixedPointTypeClass.scala 21:58]
  assign _T_47 = $signed(_T_45) + $signed(_T_39); // @[FixedPointTypeClass.scala 21:58]
  assign _T_48 = $signed(_T_47); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_8 = {{8{io_biasVecs_0_2[31]}},io_biasVecs_0_2}; // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_9 = $signed(_GEN_8) << 8; // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_10 = {{24{_GEN_9[39]}},_GEN_9}; // @[FixedPointTypeClass.scala 21:58]
  assign _T_50 = $signed(_T_48) + $signed(_GEN_10); // @[FixedPointTypeClass.scala 21:58]
  assign _T_51 = $signed(_T_50); // @[FixedPointTypeClass.scala 21:58]
  assign _T_52 = $signed(_T_51) > $signed(64'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign _T_53 = _T_52 ? $signed(_T_51) : $signed(64'sh0); // @[neuralNet.scala 50:30]
  assign _T_54 = $signed(io_in_bits_0) * $signed(io_inputWeights_3_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_55 = $signed(io_in_bits_1) * $signed(io_inputWeights_3_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_56 = $signed(io_in_bits_2) * $signed(io_inputWeights_3_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_57 = $signed(io_in_bits_3) * $signed(io_inputWeights_3_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_59 = $signed(_T_54) + $signed(_T_55); // @[FixedPointTypeClass.scala 21:58]
  assign _T_60 = $signed(_T_59); // @[FixedPointTypeClass.scala 21:58]
  assign _T_62 = $signed(_T_60) + $signed(_T_56); // @[FixedPointTypeClass.scala 21:58]
  assign _T_63 = $signed(_T_62); // @[FixedPointTypeClass.scala 21:58]
  assign _T_65 = $signed(_T_63) + $signed(_T_57); // @[FixedPointTypeClass.scala 21:58]
  assign _T_66 = $signed(_T_65); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_11 = {{8{io_biasVecs_0_3[31]}},io_biasVecs_0_3}; // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_12 = $signed(_GEN_11) << 8; // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_13 = {{24{_GEN_12[39]}},_GEN_12}; // @[FixedPointTypeClass.scala 21:58]
  assign _T_68 = $signed(_T_66) + $signed(_GEN_13); // @[FixedPointTypeClass.scala 21:58]
  assign _T_69 = $signed(_T_68); // @[FixedPointTypeClass.scala 21:58]
  assign _T_70 = $signed(_T_69) > $signed(64'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign _T_71 = _T_70 ? $signed(_T_69) : $signed(64'sh0); // @[neuralNet.scala 50:30]
  assign _T_72 = $signed(io_in_bits_0) * $signed(io_inputWeights_4_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_73 = $signed(io_in_bits_1) * $signed(io_inputWeights_4_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_74 = $signed(io_in_bits_2) * $signed(io_inputWeights_4_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_75 = $signed(io_in_bits_3) * $signed(io_inputWeights_4_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_77 = $signed(_T_72) + $signed(_T_73); // @[FixedPointTypeClass.scala 21:58]
  assign _T_78 = $signed(_T_77); // @[FixedPointTypeClass.scala 21:58]
  assign _T_80 = $signed(_T_78) + $signed(_T_74); // @[FixedPointTypeClass.scala 21:58]
  assign _T_81 = $signed(_T_80); // @[FixedPointTypeClass.scala 21:58]
  assign _T_83 = $signed(_T_81) + $signed(_T_75); // @[FixedPointTypeClass.scala 21:58]
  assign _T_84 = $signed(_T_83); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_14 = {{8{io_biasVecs_0_4[31]}},io_biasVecs_0_4}; // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_15 = $signed(_GEN_14) << 8; // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_16 = {{24{_GEN_15[39]}},_GEN_15}; // @[FixedPointTypeClass.scala 21:58]
  assign _T_86 = $signed(_T_84) + $signed(_GEN_16); // @[FixedPointTypeClass.scala 21:58]
  assign _T_87 = $signed(_T_86); // @[FixedPointTypeClass.scala 21:58]
  assign _T_88 = $signed(_T_87) > $signed(64'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign _T_89 = _T_88 ? $signed(_T_87) : $signed(64'sh0); // @[neuralNet.scala 50:30]
  assign _T_90 = $signed(io_in_bits_0) * $signed(io_inputWeights_5_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_91 = $signed(io_in_bits_1) * $signed(io_inputWeights_5_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_92 = $signed(io_in_bits_2) * $signed(io_inputWeights_5_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_93 = $signed(io_in_bits_3) * $signed(io_inputWeights_5_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_95 = $signed(_T_90) + $signed(_T_91); // @[FixedPointTypeClass.scala 21:58]
  assign _T_96 = $signed(_T_95); // @[FixedPointTypeClass.scala 21:58]
  assign _T_98 = $signed(_T_96) + $signed(_T_92); // @[FixedPointTypeClass.scala 21:58]
  assign _T_99 = $signed(_T_98); // @[FixedPointTypeClass.scala 21:58]
  assign _T_101 = $signed(_T_99) + $signed(_T_93); // @[FixedPointTypeClass.scala 21:58]
  assign _T_102 = $signed(_T_101); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_17 = {{8{io_biasVecs_0_5[31]}},io_biasVecs_0_5}; // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_18 = $signed(_GEN_17) << 8; // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_19 = {{24{_GEN_18[39]}},_GEN_18}; // @[FixedPointTypeClass.scala 21:58]
  assign _T_104 = $signed(_T_102) + $signed(_GEN_19); // @[FixedPointTypeClass.scala 21:58]
  assign _T_105 = $signed(_T_104); // @[FixedPointTypeClass.scala 21:58]
  assign _T_106 = $signed(_T_105) > $signed(64'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign _T_107 = _T_106 ? $signed(_T_105) : $signed(64'sh0); // @[neuralNet.scala 50:30]
  assign _T_108 = $signed(io_in_bits_0) * $signed(io_inputWeights_6_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_109 = $signed(io_in_bits_1) * $signed(io_inputWeights_6_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_110 = $signed(io_in_bits_2) * $signed(io_inputWeights_6_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_111 = $signed(io_in_bits_3) * $signed(io_inputWeights_6_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_113 = $signed(_T_108) + $signed(_T_109); // @[FixedPointTypeClass.scala 21:58]
  assign _T_114 = $signed(_T_113); // @[FixedPointTypeClass.scala 21:58]
  assign _T_116 = $signed(_T_114) + $signed(_T_110); // @[FixedPointTypeClass.scala 21:58]
  assign _T_117 = $signed(_T_116); // @[FixedPointTypeClass.scala 21:58]
  assign _T_119 = $signed(_T_117) + $signed(_T_111); // @[FixedPointTypeClass.scala 21:58]
  assign _T_120 = $signed(_T_119); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_20 = {{8{io_biasVecs_0_6[31]}},io_biasVecs_0_6}; // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_21 = $signed(_GEN_20) << 8; // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_22 = {{24{_GEN_21[39]}},_GEN_21}; // @[FixedPointTypeClass.scala 21:58]
  assign _T_122 = $signed(_T_120) + $signed(_GEN_22); // @[FixedPointTypeClass.scala 21:58]
  assign _T_123 = $signed(_T_122); // @[FixedPointTypeClass.scala 21:58]
  assign _T_124 = $signed(_T_123) > $signed(64'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign _T_125 = _T_124 ? $signed(_T_123) : $signed(64'sh0); // @[neuralNet.scala 50:30]
  assign _T_126 = $signed(io_in_bits_0) * $signed(io_inputWeights_7_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_127 = $signed(io_in_bits_1) * $signed(io_inputWeights_7_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_128 = $signed(io_in_bits_2) * $signed(io_inputWeights_7_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_129 = $signed(io_in_bits_3) * $signed(io_inputWeights_7_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_131 = $signed(_T_126) + $signed(_T_127); // @[FixedPointTypeClass.scala 21:58]
  assign _T_132 = $signed(_T_131); // @[FixedPointTypeClass.scala 21:58]
  assign _T_134 = $signed(_T_132) + $signed(_T_128); // @[FixedPointTypeClass.scala 21:58]
  assign _T_135 = $signed(_T_134); // @[FixedPointTypeClass.scala 21:58]
  assign _T_137 = $signed(_T_135) + $signed(_T_129); // @[FixedPointTypeClass.scala 21:58]
  assign _T_138 = $signed(_T_137); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_23 = {{8{io_biasVecs_0_7[31]}},io_biasVecs_0_7}; // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_24 = $signed(_GEN_23) << 8; // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_25 = {{24{_GEN_24[39]}},_GEN_24}; // @[FixedPointTypeClass.scala 21:58]
  assign _T_140 = $signed(_T_138) + $signed(_GEN_25); // @[FixedPointTypeClass.scala 21:58]
  assign _T_141 = $signed(_T_140); // @[FixedPointTypeClass.scala 21:58]
  assign _T_142 = $signed(_T_141) > $signed(64'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign _T_143 = _T_142 ? $signed(_T_141) : $signed(64'sh0); // @[neuralNet.scala 50:30]
  assign _T_144 = $signed(io_in_bits_0) * $signed(io_inputWeights_8_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_145 = $signed(io_in_bits_1) * $signed(io_inputWeights_8_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_146 = $signed(io_in_bits_2) * $signed(io_inputWeights_8_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_147 = $signed(io_in_bits_3) * $signed(io_inputWeights_8_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_149 = $signed(_T_144) + $signed(_T_145); // @[FixedPointTypeClass.scala 21:58]
  assign _T_150 = $signed(_T_149); // @[FixedPointTypeClass.scala 21:58]
  assign _T_152 = $signed(_T_150) + $signed(_T_146); // @[FixedPointTypeClass.scala 21:58]
  assign _T_153 = $signed(_T_152); // @[FixedPointTypeClass.scala 21:58]
  assign _T_155 = $signed(_T_153) + $signed(_T_147); // @[FixedPointTypeClass.scala 21:58]
  assign _T_156 = $signed(_T_155); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_26 = {{8{io_biasVecs_0_8[31]}},io_biasVecs_0_8}; // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_27 = $signed(_GEN_26) << 8; // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_28 = {{24{_GEN_27[39]}},_GEN_27}; // @[FixedPointTypeClass.scala 21:58]
  assign _T_158 = $signed(_T_156) + $signed(_GEN_28); // @[FixedPointTypeClass.scala 21:58]
  assign _T_159 = $signed(_T_158); // @[FixedPointTypeClass.scala 21:58]
  assign _T_160 = $signed(_T_159) > $signed(64'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign _T_161 = _T_160 ? $signed(_T_159) : $signed(64'sh0); // @[neuralNet.scala 50:30]
  assign _T_162 = $signed(io_in_bits_0) * $signed(io_inputWeights_9_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_163 = $signed(io_in_bits_1) * $signed(io_inputWeights_9_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_164 = $signed(io_in_bits_2) * $signed(io_inputWeights_9_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_165 = $signed(io_in_bits_3) * $signed(io_inputWeights_9_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_167 = $signed(_T_162) + $signed(_T_163); // @[FixedPointTypeClass.scala 21:58]
  assign _T_168 = $signed(_T_167); // @[FixedPointTypeClass.scala 21:58]
  assign _T_170 = $signed(_T_168) + $signed(_T_164); // @[FixedPointTypeClass.scala 21:58]
  assign _T_171 = $signed(_T_170); // @[FixedPointTypeClass.scala 21:58]
  assign _T_173 = $signed(_T_171) + $signed(_T_165); // @[FixedPointTypeClass.scala 21:58]
  assign _T_174 = $signed(_T_173); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_29 = {{8{io_biasVecs_0_9[31]}},io_biasVecs_0_9}; // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_30 = $signed(_GEN_29) << 8; // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_31 = {{24{_GEN_30[39]}},_GEN_30}; // @[FixedPointTypeClass.scala 21:58]
  assign _T_176 = $signed(_T_174) + $signed(_GEN_31); // @[FixedPointTypeClass.scala 21:58]
  assign _T_177 = $signed(_T_176); // @[FixedPointTypeClass.scala 21:58]
  assign _T_178 = $signed(_T_177) > $signed(64'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign _T_179 = _T_178 ? $signed(_T_177) : $signed(64'sh0); // @[neuralNet.scala 50:30]
  assign _GEN_32 = _T_17[63:8]; // @[neuralNet.scala 43:26 neuralNet.scala 50:24]
  assign _GEN_33 = _GEN_32[31:0]; // @[neuralNet.scala 43:26 neuralNet.scala 50:24]
  assign hiddenLayers_0_0 = $signed(_GEN_33); // @[neuralNet.scala 43:26 neuralNet.scala 50:24]
  assign _T_180 = $signed(hiddenLayers_0_0) * $signed(io_midAndOutputWeights_0_0); // @[FixedPointTypeClass.scala 43:59]
  assign _GEN_34 = _T_35[63:8]; // @[neuralNet.scala 43:26 neuralNet.scala 50:24]
  assign _GEN_35 = _GEN_34[31:0]; // @[neuralNet.scala 43:26 neuralNet.scala 50:24]
  assign hiddenLayers_0_1 = $signed(_GEN_35); // @[neuralNet.scala 43:26 neuralNet.scala 50:24]
  assign _T_181 = $signed(hiddenLayers_0_1) * $signed(io_midAndOutputWeights_0_1); // @[FixedPointTypeClass.scala 43:59]
  assign _GEN_36 = _T_53[63:8]; // @[neuralNet.scala 43:26 neuralNet.scala 50:24]
  assign _GEN_37 = _GEN_36[31:0]; // @[neuralNet.scala 43:26 neuralNet.scala 50:24]
  assign hiddenLayers_0_2 = $signed(_GEN_37); // @[neuralNet.scala 43:26 neuralNet.scala 50:24]
  assign _T_182 = $signed(hiddenLayers_0_2) * $signed(io_midAndOutputWeights_0_2); // @[FixedPointTypeClass.scala 43:59]
  assign _GEN_38 = _T_71[63:8]; // @[neuralNet.scala 43:26 neuralNet.scala 50:24]
  assign _GEN_39 = _GEN_38[31:0]; // @[neuralNet.scala 43:26 neuralNet.scala 50:24]
  assign hiddenLayers_0_3 = $signed(_GEN_39); // @[neuralNet.scala 43:26 neuralNet.scala 50:24]
  assign _T_183 = $signed(hiddenLayers_0_3) * $signed(io_midAndOutputWeights_0_3); // @[FixedPointTypeClass.scala 43:59]
  assign _GEN_40 = _T_89[63:8]; // @[neuralNet.scala 43:26 neuralNet.scala 50:24]
  assign _GEN_41 = _GEN_40[31:0]; // @[neuralNet.scala 43:26 neuralNet.scala 50:24]
  assign hiddenLayers_0_4 = $signed(_GEN_41); // @[neuralNet.scala 43:26 neuralNet.scala 50:24]
  assign _T_184 = $signed(hiddenLayers_0_4) * $signed(io_midAndOutputWeights_0_4); // @[FixedPointTypeClass.scala 43:59]
  assign _GEN_42 = _T_107[63:8]; // @[neuralNet.scala 43:26 neuralNet.scala 50:24]
  assign _GEN_43 = _GEN_42[31:0]; // @[neuralNet.scala 43:26 neuralNet.scala 50:24]
  assign hiddenLayers_0_5 = $signed(_GEN_43); // @[neuralNet.scala 43:26 neuralNet.scala 50:24]
  assign _T_185 = $signed(hiddenLayers_0_5) * $signed(io_midAndOutputWeights_0_5); // @[FixedPointTypeClass.scala 43:59]
  assign _GEN_44 = _T_125[63:8]; // @[neuralNet.scala 43:26 neuralNet.scala 50:24]
  assign _GEN_45 = _GEN_44[31:0]; // @[neuralNet.scala 43:26 neuralNet.scala 50:24]
  assign hiddenLayers_0_6 = $signed(_GEN_45); // @[neuralNet.scala 43:26 neuralNet.scala 50:24]
  assign _T_186 = $signed(hiddenLayers_0_6) * $signed(io_midAndOutputWeights_0_6); // @[FixedPointTypeClass.scala 43:59]
  assign _GEN_46 = _T_143[63:8]; // @[neuralNet.scala 43:26 neuralNet.scala 50:24]
  assign _GEN_47 = _GEN_46[31:0]; // @[neuralNet.scala 43:26 neuralNet.scala 50:24]
  assign hiddenLayers_0_7 = $signed(_GEN_47); // @[neuralNet.scala 43:26 neuralNet.scala 50:24]
  assign _T_187 = $signed(hiddenLayers_0_7) * $signed(io_midAndOutputWeights_0_7); // @[FixedPointTypeClass.scala 43:59]
  assign _GEN_48 = _T_161[63:8]; // @[neuralNet.scala 43:26 neuralNet.scala 50:24]
  assign _GEN_49 = _GEN_48[31:0]; // @[neuralNet.scala 43:26 neuralNet.scala 50:24]
  assign hiddenLayers_0_8 = $signed(_GEN_49); // @[neuralNet.scala 43:26 neuralNet.scala 50:24]
  assign _T_188 = $signed(hiddenLayers_0_8) * $signed(io_midAndOutputWeights_0_8); // @[FixedPointTypeClass.scala 43:59]
  assign _GEN_50 = _T_179[63:8]; // @[neuralNet.scala 43:26 neuralNet.scala 50:24]
  assign _GEN_51 = _GEN_50[31:0]; // @[neuralNet.scala 43:26 neuralNet.scala 50:24]
  assign hiddenLayers_0_9 = $signed(_GEN_51); // @[neuralNet.scala 43:26 neuralNet.scala 50:24]
  assign _T_189 = $signed(hiddenLayers_0_9) * $signed(io_midAndOutputWeights_0_9); // @[FixedPointTypeClass.scala 43:59]
  assign _T_191 = $signed(_T_180) + $signed(_T_181); // @[FixedPointTypeClass.scala 21:58]
  assign _T_192 = $signed(_T_191); // @[FixedPointTypeClass.scala 21:58]
  assign _T_194 = $signed(_T_192) + $signed(_T_182); // @[FixedPointTypeClass.scala 21:58]
  assign _T_195 = $signed(_T_194); // @[FixedPointTypeClass.scala 21:58]
  assign _T_197 = $signed(_T_195) + $signed(_T_183); // @[FixedPointTypeClass.scala 21:58]
  assign _T_198 = $signed(_T_197); // @[FixedPointTypeClass.scala 21:58]
  assign _T_200 = $signed(_T_198) + $signed(_T_184); // @[FixedPointTypeClass.scala 21:58]
  assign _T_201 = $signed(_T_200); // @[FixedPointTypeClass.scala 21:58]
  assign _T_203 = $signed(_T_201) + $signed(_T_185); // @[FixedPointTypeClass.scala 21:58]
  assign _T_204 = $signed(_T_203); // @[FixedPointTypeClass.scala 21:58]
  assign _T_206 = $signed(_T_204) + $signed(_T_186); // @[FixedPointTypeClass.scala 21:58]
  assign _T_207 = $signed(_T_206); // @[FixedPointTypeClass.scala 21:58]
  assign _T_209 = $signed(_T_207) + $signed(_T_187); // @[FixedPointTypeClass.scala 21:58]
  assign _T_210 = $signed(_T_209); // @[FixedPointTypeClass.scala 21:58]
  assign _T_212 = $signed(_T_210) + $signed(_T_188); // @[FixedPointTypeClass.scala 21:58]
  assign _T_213 = $signed(_T_212); // @[FixedPointTypeClass.scala 21:58]
  assign _T_215 = $signed(_T_213) + $signed(_T_189); // @[FixedPointTypeClass.scala 21:58]
  assign _T_216 = $signed(_T_215); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_52 = {{8{io_biasVecs_1_0[31]}},io_biasVecs_1_0}; // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_53 = $signed(_GEN_52) << 8; // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_54 = {{24{_GEN_53[39]}},_GEN_53}; // @[FixedPointTypeClass.scala 21:58]
  assign _T_218 = $signed(_T_216) + $signed(_GEN_54); // @[FixedPointTypeClass.scala 21:58]
  assign _T_219 = $signed(_T_218); // @[FixedPointTypeClass.scala 21:58]
  assign _T_220 = $signed(_T_219) > $signed(64'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign _T_221 = _T_220 ? $signed(_T_219) : $signed(64'sh0); // @[neuralNet.scala 59:32]
  assign _T_222 = $signed(hiddenLayers_0_0) * $signed(io_midAndOutputWeights_1_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_223 = $signed(hiddenLayers_0_1) * $signed(io_midAndOutputWeights_1_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_224 = $signed(hiddenLayers_0_2) * $signed(io_midAndOutputWeights_1_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_225 = $signed(hiddenLayers_0_3) * $signed(io_midAndOutputWeights_1_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_226 = $signed(hiddenLayers_0_4) * $signed(io_midAndOutputWeights_1_4); // @[FixedPointTypeClass.scala 43:59]
  assign _T_227 = $signed(hiddenLayers_0_5) * $signed(io_midAndOutputWeights_1_5); // @[FixedPointTypeClass.scala 43:59]
  assign _T_228 = $signed(hiddenLayers_0_6) * $signed(io_midAndOutputWeights_1_6); // @[FixedPointTypeClass.scala 43:59]
  assign _T_229 = $signed(hiddenLayers_0_7) * $signed(io_midAndOutputWeights_1_7); // @[FixedPointTypeClass.scala 43:59]
  assign _T_230 = $signed(hiddenLayers_0_8) * $signed(io_midAndOutputWeights_1_8); // @[FixedPointTypeClass.scala 43:59]
  assign _T_231 = $signed(hiddenLayers_0_9) * $signed(io_midAndOutputWeights_1_9); // @[FixedPointTypeClass.scala 43:59]
  assign _T_233 = $signed(_T_222) + $signed(_T_223); // @[FixedPointTypeClass.scala 21:58]
  assign _T_234 = $signed(_T_233); // @[FixedPointTypeClass.scala 21:58]
  assign _T_236 = $signed(_T_234) + $signed(_T_224); // @[FixedPointTypeClass.scala 21:58]
  assign _T_237 = $signed(_T_236); // @[FixedPointTypeClass.scala 21:58]
  assign _T_239 = $signed(_T_237) + $signed(_T_225); // @[FixedPointTypeClass.scala 21:58]
  assign _T_240 = $signed(_T_239); // @[FixedPointTypeClass.scala 21:58]
  assign _T_242 = $signed(_T_240) + $signed(_T_226); // @[FixedPointTypeClass.scala 21:58]
  assign _T_243 = $signed(_T_242); // @[FixedPointTypeClass.scala 21:58]
  assign _T_245 = $signed(_T_243) + $signed(_T_227); // @[FixedPointTypeClass.scala 21:58]
  assign _T_246 = $signed(_T_245); // @[FixedPointTypeClass.scala 21:58]
  assign _T_248 = $signed(_T_246) + $signed(_T_228); // @[FixedPointTypeClass.scala 21:58]
  assign _T_249 = $signed(_T_248); // @[FixedPointTypeClass.scala 21:58]
  assign _T_251 = $signed(_T_249) + $signed(_T_229); // @[FixedPointTypeClass.scala 21:58]
  assign _T_252 = $signed(_T_251); // @[FixedPointTypeClass.scala 21:58]
  assign _T_254 = $signed(_T_252) + $signed(_T_230); // @[FixedPointTypeClass.scala 21:58]
  assign _T_255 = $signed(_T_254); // @[FixedPointTypeClass.scala 21:58]
  assign _T_257 = $signed(_T_255) + $signed(_T_231); // @[FixedPointTypeClass.scala 21:58]
  assign _T_258 = $signed(_T_257); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_55 = {{8{io_biasVecs_1_1[31]}},io_biasVecs_1_1}; // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_56 = $signed(_GEN_55) << 8; // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_57 = {{24{_GEN_56[39]}},_GEN_56}; // @[FixedPointTypeClass.scala 21:58]
  assign _T_260 = $signed(_T_258) + $signed(_GEN_57); // @[FixedPointTypeClass.scala 21:58]
  assign _T_261 = $signed(_T_260); // @[FixedPointTypeClass.scala 21:58]
  assign _T_262 = $signed(_T_261) > $signed(64'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign _T_263 = _T_262 ? $signed(_T_261) : $signed(64'sh0); // @[neuralNet.scala 59:32]
  assign _T_264 = $signed(hiddenLayers_0_0) * $signed(io_midAndOutputWeights_2_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_265 = $signed(hiddenLayers_0_1) * $signed(io_midAndOutputWeights_2_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_266 = $signed(hiddenLayers_0_2) * $signed(io_midAndOutputWeights_2_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_267 = $signed(hiddenLayers_0_3) * $signed(io_midAndOutputWeights_2_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_268 = $signed(hiddenLayers_0_4) * $signed(io_midAndOutputWeights_2_4); // @[FixedPointTypeClass.scala 43:59]
  assign _T_269 = $signed(hiddenLayers_0_5) * $signed(io_midAndOutputWeights_2_5); // @[FixedPointTypeClass.scala 43:59]
  assign _T_270 = $signed(hiddenLayers_0_6) * $signed(io_midAndOutputWeights_2_6); // @[FixedPointTypeClass.scala 43:59]
  assign _T_271 = $signed(hiddenLayers_0_7) * $signed(io_midAndOutputWeights_2_7); // @[FixedPointTypeClass.scala 43:59]
  assign _T_272 = $signed(hiddenLayers_0_8) * $signed(io_midAndOutputWeights_2_8); // @[FixedPointTypeClass.scala 43:59]
  assign _T_273 = $signed(hiddenLayers_0_9) * $signed(io_midAndOutputWeights_2_9); // @[FixedPointTypeClass.scala 43:59]
  assign _T_275 = $signed(_T_264) + $signed(_T_265); // @[FixedPointTypeClass.scala 21:58]
  assign _T_276 = $signed(_T_275); // @[FixedPointTypeClass.scala 21:58]
  assign _T_278 = $signed(_T_276) + $signed(_T_266); // @[FixedPointTypeClass.scala 21:58]
  assign _T_279 = $signed(_T_278); // @[FixedPointTypeClass.scala 21:58]
  assign _T_281 = $signed(_T_279) + $signed(_T_267); // @[FixedPointTypeClass.scala 21:58]
  assign _T_282 = $signed(_T_281); // @[FixedPointTypeClass.scala 21:58]
  assign _T_284 = $signed(_T_282) + $signed(_T_268); // @[FixedPointTypeClass.scala 21:58]
  assign _T_285 = $signed(_T_284); // @[FixedPointTypeClass.scala 21:58]
  assign _T_287 = $signed(_T_285) + $signed(_T_269); // @[FixedPointTypeClass.scala 21:58]
  assign _T_288 = $signed(_T_287); // @[FixedPointTypeClass.scala 21:58]
  assign _T_290 = $signed(_T_288) + $signed(_T_270); // @[FixedPointTypeClass.scala 21:58]
  assign _T_291 = $signed(_T_290); // @[FixedPointTypeClass.scala 21:58]
  assign _T_293 = $signed(_T_291) + $signed(_T_271); // @[FixedPointTypeClass.scala 21:58]
  assign _T_294 = $signed(_T_293); // @[FixedPointTypeClass.scala 21:58]
  assign _T_296 = $signed(_T_294) + $signed(_T_272); // @[FixedPointTypeClass.scala 21:58]
  assign _T_297 = $signed(_T_296); // @[FixedPointTypeClass.scala 21:58]
  assign _T_299 = $signed(_T_297) + $signed(_T_273); // @[FixedPointTypeClass.scala 21:58]
  assign _T_300 = $signed(_T_299); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_58 = {{8{io_biasVecs_1_2[31]}},io_biasVecs_1_2}; // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_59 = $signed(_GEN_58) << 8; // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_60 = {{24{_GEN_59[39]}},_GEN_59}; // @[FixedPointTypeClass.scala 21:58]
  assign _T_302 = $signed(_T_300) + $signed(_GEN_60); // @[FixedPointTypeClass.scala 21:58]
  assign _T_303 = $signed(_T_302); // @[FixedPointTypeClass.scala 21:58]
  assign _T_304 = $signed(_T_303) > $signed(64'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign _T_305 = _T_304 ? $signed(_T_303) : $signed(64'sh0); // @[neuralNet.scala 59:32]
  assign _T_306 = $signed(hiddenLayers_0_0) * $signed(io_midAndOutputWeights_3_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_307 = $signed(hiddenLayers_0_1) * $signed(io_midAndOutputWeights_3_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_308 = $signed(hiddenLayers_0_2) * $signed(io_midAndOutputWeights_3_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_309 = $signed(hiddenLayers_0_3) * $signed(io_midAndOutputWeights_3_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_310 = $signed(hiddenLayers_0_4) * $signed(io_midAndOutputWeights_3_4); // @[FixedPointTypeClass.scala 43:59]
  assign _T_311 = $signed(hiddenLayers_0_5) * $signed(io_midAndOutputWeights_3_5); // @[FixedPointTypeClass.scala 43:59]
  assign _T_312 = $signed(hiddenLayers_0_6) * $signed(io_midAndOutputWeights_3_6); // @[FixedPointTypeClass.scala 43:59]
  assign _T_313 = $signed(hiddenLayers_0_7) * $signed(io_midAndOutputWeights_3_7); // @[FixedPointTypeClass.scala 43:59]
  assign _T_314 = $signed(hiddenLayers_0_8) * $signed(io_midAndOutputWeights_3_8); // @[FixedPointTypeClass.scala 43:59]
  assign _T_315 = $signed(hiddenLayers_0_9) * $signed(io_midAndOutputWeights_3_9); // @[FixedPointTypeClass.scala 43:59]
  assign _T_317 = $signed(_T_306) + $signed(_T_307); // @[FixedPointTypeClass.scala 21:58]
  assign _T_318 = $signed(_T_317); // @[FixedPointTypeClass.scala 21:58]
  assign _T_320 = $signed(_T_318) + $signed(_T_308); // @[FixedPointTypeClass.scala 21:58]
  assign _T_321 = $signed(_T_320); // @[FixedPointTypeClass.scala 21:58]
  assign _T_323 = $signed(_T_321) + $signed(_T_309); // @[FixedPointTypeClass.scala 21:58]
  assign _T_324 = $signed(_T_323); // @[FixedPointTypeClass.scala 21:58]
  assign _T_326 = $signed(_T_324) + $signed(_T_310); // @[FixedPointTypeClass.scala 21:58]
  assign _T_327 = $signed(_T_326); // @[FixedPointTypeClass.scala 21:58]
  assign _T_329 = $signed(_T_327) + $signed(_T_311); // @[FixedPointTypeClass.scala 21:58]
  assign _T_330 = $signed(_T_329); // @[FixedPointTypeClass.scala 21:58]
  assign _T_332 = $signed(_T_330) + $signed(_T_312); // @[FixedPointTypeClass.scala 21:58]
  assign _T_333 = $signed(_T_332); // @[FixedPointTypeClass.scala 21:58]
  assign _T_335 = $signed(_T_333) + $signed(_T_313); // @[FixedPointTypeClass.scala 21:58]
  assign _T_336 = $signed(_T_335); // @[FixedPointTypeClass.scala 21:58]
  assign _T_338 = $signed(_T_336) + $signed(_T_314); // @[FixedPointTypeClass.scala 21:58]
  assign _T_339 = $signed(_T_338); // @[FixedPointTypeClass.scala 21:58]
  assign _T_341 = $signed(_T_339) + $signed(_T_315); // @[FixedPointTypeClass.scala 21:58]
  assign _T_342 = $signed(_T_341); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_61 = {{8{io_biasVecs_1_3[31]}},io_biasVecs_1_3}; // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_62 = $signed(_GEN_61) << 8; // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_63 = {{24{_GEN_62[39]}},_GEN_62}; // @[FixedPointTypeClass.scala 21:58]
  assign _T_344 = $signed(_T_342) + $signed(_GEN_63); // @[FixedPointTypeClass.scala 21:58]
  assign _T_345 = $signed(_T_344); // @[FixedPointTypeClass.scala 21:58]
  assign _T_346 = $signed(_T_345) > $signed(64'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign _T_347 = _T_346 ? $signed(_T_345) : $signed(64'sh0); // @[neuralNet.scala 59:32]
  assign _T_348 = $signed(hiddenLayers_0_0) * $signed(io_midAndOutputWeights_4_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_349 = $signed(hiddenLayers_0_1) * $signed(io_midAndOutputWeights_4_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_350 = $signed(hiddenLayers_0_2) * $signed(io_midAndOutputWeights_4_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_351 = $signed(hiddenLayers_0_3) * $signed(io_midAndOutputWeights_4_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_352 = $signed(hiddenLayers_0_4) * $signed(io_midAndOutputWeights_4_4); // @[FixedPointTypeClass.scala 43:59]
  assign _T_353 = $signed(hiddenLayers_0_5) * $signed(io_midAndOutputWeights_4_5); // @[FixedPointTypeClass.scala 43:59]
  assign _T_354 = $signed(hiddenLayers_0_6) * $signed(io_midAndOutputWeights_4_6); // @[FixedPointTypeClass.scala 43:59]
  assign _T_355 = $signed(hiddenLayers_0_7) * $signed(io_midAndOutputWeights_4_7); // @[FixedPointTypeClass.scala 43:59]
  assign _T_356 = $signed(hiddenLayers_0_8) * $signed(io_midAndOutputWeights_4_8); // @[FixedPointTypeClass.scala 43:59]
  assign _T_357 = $signed(hiddenLayers_0_9) * $signed(io_midAndOutputWeights_4_9); // @[FixedPointTypeClass.scala 43:59]
  assign _T_359 = $signed(_T_348) + $signed(_T_349); // @[FixedPointTypeClass.scala 21:58]
  assign _T_360 = $signed(_T_359); // @[FixedPointTypeClass.scala 21:58]
  assign _T_362 = $signed(_T_360) + $signed(_T_350); // @[FixedPointTypeClass.scala 21:58]
  assign _T_363 = $signed(_T_362); // @[FixedPointTypeClass.scala 21:58]
  assign _T_365 = $signed(_T_363) + $signed(_T_351); // @[FixedPointTypeClass.scala 21:58]
  assign _T_366 = $signed(_T_365); // @[FixedPointTypeClass.scala 21:58]
  assign _T_368 = $signed(_T_366) + $signed(_T_352); // @[FixedPointTypeClass.scala 21:58]
  assign _T_369 = $signed(_T_368); // @[FixedPointTypeClass.scala 21:58]
  assign _T_371 = $signed(_T_369) + $signed(_T_353); // @[FixedPointTypeClass.scala 21:58]
  assign _T_372 = $signed(_T_371); // @[FixedPointTypeClass.scala 21:58]
  assign _T_374 = $signed(_T_372) + $signed(_T_354); // @[FixedPointTypeClass.scala 21:58]
  assign _T_375 = $signed(_T_374); // @[FixedPointTypeClass.scala 21:58]
  assign _T_377 = $signed(_T_375) + $signed(_T_355); // @[FixedPointTypeClass.scala 21:58]
  assign _T_378 = $signed(_T_377); // @[FixedPointTypeClass.scala 21:58]
  assign _T_380 = $signed(_T_378) + $signed(_T_356); // @[FixedPointTypeClass.scala 21:58]
  assign _T_381 = $signed(_T_380); // @[FixedPointTypeClass.scala 21:58]
  assign _T_383 = $signed(_T_381) + $signed(_T_357); // @[FixedPointTypeClass.scala 21:58]
  assign _T_384 = $signed(_T_383); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_64 = {{8{io_biasVecs_1_4[31]}},io_biasVecs_1_4}; // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_65 = $signed(_GEN_64) << 8; // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_66 = {{24{_GEN_65[39]}},_GEN_65}; // @[FixedPointTypeClass.scala 21:58]
  assign _T_386 = $signed(_T_384) + $signed(_GEN_66); // @[FixedPointTypeClass.scala 21:58]
  assign _T_387 = $signed(_T_386); // @[FixedPointTypeClass.scala 21:58]
  assign _T_388 = $signed(_T_387) > $signed(64'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign _T_389 = _T_388 ? $signed(_T_387) : $signed(64'sh0); // @[neuralNet.scala 59:32]
  assign _T_390 = $signed(hiddenLayers_0_0) * $signed(io_midAndOutputWeights_5_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_391 = $signed(hiddenLayers_0_1) * $signed(io_midAndOutputWeights_5_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_392 = $signed(hiddenLayers_0_2) * $signed(io_midAndOutputWeights_5_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_393 = $signed(hiddenLayers_0_3) * $signed(io_midAndOutputWeights_5_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_394 = $signed(hiddenLayers_0_4) * $signed(io_midAndOutputWeights_5_4); // @[FixedPointTypeClass.scala 43:59]
  assign _T_395 = $signed(hiddenLayers_0_5) * $signed(io_midAndOutputWeights_5_5); // @[FixedPointTypeClass.scala 43:59]
  assign _T_396 = $signed(hiddenLayers_0_6) * $signed(io_midAndOutputWeights_5_6); // @[FixedPointTypeClass.scala 43:59]
  assign _T_397 = $signed(hiddenLayers_0_7) * $signed(io_midAndOutputWeights_5_7); // @[FixedPointTypeClass.scala 43:59]
  assign _T_398 = $signed(hiddenLayers_0_8) * $signed(io_midAndOutputWeights_5_8); // @[FixedPointTypeClass.scala 43:59]
  assign _T_399 = $signed(hiddenLayers_0_9) * $signed(io_midAndOutputWeights_5_9); // @[FixedPointTypeClass.scala 43:59]
  assign _T_401 = $signed(_T_390) + $signed(_T_391); // @[FixedPointTypeClass.scala 21:58]
  assign _T_402 = $signed(_T_401); // @[FixedPointTypeClass.scala 21:58]
  assign _T_404 = $signed(_T_402) + $signed(_T_392); // @[FixedPointTypeClass.scala 21:58]
  assign _T_405 = $signed(_T_404); // @[FixedPointTypeClass.scala 21:58]
  assign _T_407 = $signed(_T_405) + $signed(_T_393); // @[FixedPointTypeClass.scala 21:58]
  assign _T_408 = $signed(_T_407); // @[FixedPointTypeClass.scala 21:58]
  assign _T_410 = $signed(_T_408) + $signed(_T_394); // @[FixedPointTypeClass.scala 21:58]
  assign _T_411 = $signed(_T_410); // @[FixedPointTypeClass.scala 21:58]
  assign _T_413 = $signed(_T_411) + $signed(_T_395); // @[FixedPointTypeClass.scala 21:58]
  assign _T_414 = $signed(_T_413); // @[FixedPointTypeClass.scala 21:58]
  assign _T_416 = $signed(_T_414) + $signed(_T_396); // @[FixedPointTypeClass.scala 21:58]
  assign _T_417 = $signed(_T_416); // @[FixedPointTypeClass.scala 21:58]
  assign _T_419 = $signed(_T_417) + $signed(_T_397); // @[FixedPointTypeClass.scala 21:58]
  assign _T_420 = $signed(_T_419); // @[FixedPointTypeClass.scala 21:58]
  assign _T_422 = $signed(_T_420) + $signed(_T_398); // @[FixedPointTypeClass.scala 21:58]
  assign _T_423 = $signed(_T_422); // @[FixedPointTypeClass.scala 21:58]
  assign _T_425 = $signed(_T_423) + $signed(_T_399); // @[FixedPointTypeClass.scala 21:58]
  assign _T_426 = $signed(_T_425); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_67 = {{8{io_biasVecs_1_5[31]}},io_biasVecs_1_5}; // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_68 = $signed(_GEN_67) << 8; // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_69 = {{24{_GEN_68[39]}},_GEN_68}; // @[FixedPointTypeClass.scala 21:58]
  assign _T_428 = $signed(_T_426) + $signed(_GEN_69); // @[FixedPointTypeClass.scala 21:58]
  assign _T_429 = $signed(_T_428); // @[FixedPointTypeClass.scala 21:58]
  assign _T_430 = $signed(_T_429) > $signed(64'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign _T_431 = _T_430 ? $signed(_T_429) : $signed(64'sh0); // @[neuralNet.scala 59:32]
  assign _T_432 = $signed(hiddenLayers_0_0) * $signed(io_midAndOutputWeights_6_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_433 = $signed(hiddenLayers_0_1) * $signed(io_midAndOutputWeights_6_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_434 = $signed(hiddenLayers_0_2) * $signed(io_midAndOutputWeights_6_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_435 = $signed(hiddenLayers_0_3) * $signed(io_midAndOutputWeights_6_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_436 = $signed(hiddenLayers_0_4) * $signed(io_midAndOutputWeights_6_4); // @[FixedPointTypeClass.scala 43:59]
  assign _T_437 = $signed(hiddenLayers_0_5) * $signed(io_midAndOutputWeights_6_5); // @[FixedPointTypeClass.scala 43:59]
  assign _T_438 = $signed(hiddenLayers_0_6) * $signed(io_midAndOutputWeights_6_6); // @[FixedPointTypeClass.scala 43:59]
  assign _T_439 = $signed(hiddenLayers_0_7) * $signed(io_midAndOutputWeights_6_7); // @[FixedPointTypeClass.scala 43:59]
  assign _T_440 = $signed(hiddenLayers_0_8) * $signed(io_midAndOutputWeights_6_8); // @[FixedPointTypeClass.scala 43:59]
  assign _T_441 = $signed(hiddenLayers_0_9) * $signed(io_midAndOutputWeights_6_9); // @[FixedPointTypeClass.scala 43:59]
  assign _T_443 = $signed(_T_432) + $signed(_T_433); // @[FixedPointTypeClass.scala 21:58]
  assign _T_444 = $signed(_T_443); // @[FixedPointTypeClass.scala 21:58]
  assign _T_446 = $signed(_T_444) + $signed(_T_434); // @[FixedPointTypeClass.scala 21:58]
  assign _T_447 = $signed(_T_446); // @[FixedPointTypeClass.scala 21:58]
  assign _T_449 = $signed(_T_447) + $signed(_T_435); // @[FixedPointTypeClass.scala 21:58]
  assign _T_450 = $signed(_T_449); // @[FixedPointTypeClass.scala 21:58]
  assign _T_452 = $signed(_T_450) + $signed(_T_436); // @[FixedPointTypeClass.scala 21:58]
  assign _T_453 = $signed(_T_452); // @[FixedPointTypeClass.scala 21:58]
  assign _T_455 = $signed(_T_453) + $signed(_T_437); // @[FixedPointTypeClass.scala 21:58]
  assign _T_456 = $signed(_T_455); // @[FixedPointTypeClass.scala 21:58]
  assign _T_458 = $signed(_T_456) + $signed(_T_438); // @[FixedPointTypeClass.scala 21:58]
  assign _T_459 = $signed(_T_458); // @[FixedPointTypeClass.scala 21:58]
  assign _T_461 = $signed(_T_459) + $signed(_T_439); // @[FixedPointTypeClass.scala 21:58]
  assign _T_462 = $signed(_T_461); // @[FixedPointTypeClass.scala 21:58]
  assign _T_464 = $signed(_T_462) + $signed(_T_440); // @[FixedPointTypeClass.scala 21:58]
  assign _T_465 = $signed(_T_464); // @[FixedPointTypeClass.scala 21:58]
  assign _T_467 = $signed(_T_465) + $signed(_T_441); // @[FixedPointTypeClass.scala 21:58]
  assign _T_468 = $signed(_T_467); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_70 = {{8{io_biasVecs_1_6[31]}},io_biasVecs_1_6}; // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_71 = $signed(_GEN_70) << 8; // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_72 = {{24{_GEN_71[39]}},_GEN_71}; // @[FixedPointTypeClass.scala 21:58]
  assign _T_470 = $signed(_T_468) + $signed(_GEN_72); // @[FixedPointTypeClass.scala 21:58]
  assign _T_471 = $signed(_T_470); // @[FixedPointTypeClass.scala 21:58]
  assign _T_472 = $signed(_T_471) > $signed(64'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign _T_473 = _T_472 ? $signed(_T_471) : $signed(64'sh0); // @[neuralNet.scala 59:32]
  assign _T_474 = $signed(hiddenLayers_0_0) * $signed(io_midAndOutputWeights_7_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_475 = $signed(hiddenLayers_0_1) * $signed(io_midAndOutputWeights_7_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_476 = $signed(hiddenLayers_0_2) * $signed(io_midAndOutputWeights_7_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_477 = $signed(hiddenLayers_0_3) * $signed(io_midAndOutputWeights_7_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_478 = $signed(hiddenLayers_0_4) * $signed(io_midAndOutputWeights_7_4); // @[FixedPointTypeClass.scala 43:59]
  assign _T_479 = $signed(hiddenLayers_0_5) * $signed(io_midAndOutputWeights_7_5); // @[FixedPointTypeClass.scala 43:59]
  assign _T_480 = $signed(hiddenLayers_0_6) * $signed(io_midAndOutputWeights_7_6); // @[FixedPointTypeClass.scala 43:59]
  assign _T_481 = $signed(hiddenLayers_0_7) * $signed(io_midAndOutputWeights_7_7); // @[FixedPointTypeClass.scala 43:59]
  assign _T_482 = $signed(hiddenLayers_0_8) * $signed(io_midAndOutputWeights_7_8); // @[FixedPointTypeClass.scala 43:59]
  assign _T_483 = $signed(hiddenLayers_0_9) * $signed(io_midAndOutputWeights_7_9); // @[FixedPointTypeClass.scala 43:59]
  assign _T_485 = $signed(_T_474) + $signed(_T_475); // @[FixedPointTypeClass.scala 21:58]
  assign _T_486 = $signed(_T_485); // @[FixedPointTypeClass.scala 21:58]
  assign _T_488 = $signed(_T_486) + $signed(_T_476); // @[FixedPointTypeClass.scala 21:58]
  assign _T_489 = $signed(_T_488); // @[FixedPointTypeClass.scala 21:58]
  assign _T_491 = $signed(_T_489) + $signed(_T_477); // @[FixedPointTypeClass.scala 21:58]
  assign _T_492 = $signed(_T_491); // @[FixedPointTypeClass.scala 21:58]
  assign _T_494 = $signed(_T_492) + $signed(_T_478); // @[FixedPointTypeClass.scala 21:58]
  assign _T_495 = $signed(_T_494); // @[FixedPointTypeClass.scala 21:58]
  assign _T_497 = $signed(_T_495) + $signed(_T_479); // @[FixedPointTypeClass.scala 21:58]
  assign _T_498 = $signed(_T_497); // @[FixedPointTypeClass.scala 21:58]
  assign _T_500 = $signed(_T_498) + $signed(_T_480); // @[FixedPointTypeClass.scala 21:58]
  assign _T_501 = $signed(_T_500); // @[FixedPointTypeClass.scala 21:58]
  assign _T_503 = $signed(_T_501) + $signed(_T_481); // @[FixedPointTypeClass.scala 21:58]
  assign _T_504 = $signed(_T_503); // @[FixedPointTypeClass.scala 21:58]
  assign _T_506 = $signed(_T_504) + $signed(_T_482); // @[FixedPointTypeClass.scala 21:58]
  assign _T_507 = $signed(_T_506); // @[FixedPointTypeClass.scala 21:58]
  assign _T_509 = $signed(_T_507) + $signed(_T_483); // @[FixedPointTypeClass.scala 21:58]
  assign _T_510 = $signed(_T_509); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_73 = {{8{io_biasVecs_1_7[31]}},io_biasVecs_1_7}; // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_74 = $signed(_GEN_73) << 8; // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_75 = {{24{_GEN_74[39]}},_GEN_74}; // @[FixedPointTypeClass.scala 21:58]
  assign _T_512 = $signed(_T_510) + $signed(_GEN_75); // @[FixedPointTypeClass.scala 21:58]
  assign _T_513 = $signed(_T_512); // @[FixedPointTypeClass.scala 21:58]
  assign _T_514 = $signed(_T_513) > $signed(64'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign _T_515 = _T_514 ? $signed(_T_513) : $signed(64'sh0); // @[neuralNet.scala 59:32]
  assign _T_516 = $signed(hiddenLayers_0_0) * $signed(io_midAndOutputWeights_8_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_517 = $signed(hiddenLayers_0_1) * $signed(io_midAndOutputWeights_8_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_518 = $signed(hiddenLayers_0_2) * $signed(io_midAndOutputWeights_8_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_519 = $signed(hiddenLayers_0_3) * $signed(io_midAndOutputWeights_8_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_520 = $signed(hiddenLayers_0_4) * $signed(io_midAndOutputWeights_8_4); // @[FixedPointTypeClass.scala 43:59]
  assign _T_521 = $signed(hiddenLayers_0_5) * $signed(io_midAndOutputWeights_8_5); // @[FixedPointTypeClass.scala 43:59]
  assign _T_522 = $signed(hiddenLayers_0_6) * $signed(io_midAndOutputWeights_8_6); // @[FixedPointTypeClass.scala 43:59]
  assign _T_523 = $signed(hiddenLayers_0_7) * $signed(io_midAndOutputWeights_8_7); // @[FixedPointTypeClass.scala 43:59]
  assign _T_524 = $signed(hiddenLayers_0_8) * $signed(io_midAndOutputWeights_8_8); // @[FixedPointTypeClass.scala 43:59]
  assign _T_525 = $signed(hiddenLayers_0_9) * $signed(io_midAndOutputWeights_8_9); // @[FixedPointTypeClass.scala 43:59]
  assign _T_527 = $signed(_T_516) + $signed(_T_517); // @[FixedPointTypeClass.scala 21:58]
  assign _T_528 = $signed(_T_527); // @[FixedPointTypeClass.scala 21:58]
  assign _T_530 = $signed(_T_528) + $signed(_T_518); // @[FixedPointTypeClass.scala 21:58]
  assign _T_531 = $signed(_T_530); // @[FixedPointTypeClass.scala 21:58]
  assign _T_533 = $signed(_T_531) + $signed(_T_519); // @[FixedPointTypeClass.scala 21:58]
  assign _T_534 = $signed(_T_533); // @[FixedPointTypeClass.scala 21:58]
  assign _T_536 = $signed(_T_534) + $signed(_T_520); // @[FixedPointTypeClass.scala 21:58]
  assign _T_537 = $signed(_T_536); // @[FixedPointTypeClass.scala 21:58]
  assign _T_539 = $signed(_T_537) + $signed(_T_521); // @[FixedPointTypeClass.scala 21:58]
  assign _T_540 = $signed(_T_539); // @[FixedPointTypeClass.scala 21:58]
  assign _T_542 = $signed(_T_540) + $signed(_T_522); // @[FixedPointTypeClass.scala 21:58]
  assign _T_543 = $signed(_T_542); // @[FixedPointTypeClass.scala 21:58]
  assign _T_545 = $signed(_T_543) + $signed(_T_523); // @[FixedPointTypeClass.scala 21:58]
  assign _T_546 = $signed(_T_545); // @[FixedPointTypeClass.scala 21:58]
  assign _T_548 = $signed(_T_546) + $signed(_T_524); // @[FixedPointTypeClass.scala 21:58]
  assign _T_549 = $signed(_T_548); // @[FixedPointTypeClass.scala 21:58]
  assign _T_551 = $signed(_T_549) + $signed(_T_525); // @[FixedPointTypeClass.scala 21:58]
  assign _T_552 = $signed(_T_551); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_76 = {{8{io_biasVecs_1_8[31]}},io_biasVecs_1_8}; // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_77 = $signed(_GEN_76) << 8; // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_78 = {{24{_GEN_77[39]}},_GEN_77}; // @[FixedPointTypeClass.scala 21:58]
  assign _T_554 = $signed(_T_552) + $signed(_GEN_78); // @[FixedPointTypeClass.scala 21:58]
  assign _T_555 = $signed(_T_554); // @[FixedPointTypeClass.scala 21:58]
  assign _T_556 = $signed(_T_555) > $signed(64'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign _T_557 = _T_556 ? $signed(_T_555) : $signed(64'sh0); // @[neuralNet.scala 59:32]
  assign _T_558 = $signed(hiddenLayers_0_0) * $signed(io_midAndOutputWeights_9_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_559 = $signed(hiddenLayers_0_1) * $signed(io_midAndOutputWeights_9_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_560 = $signed(hiddenLayers_0_2) * $signed(io_midAndOutputWeights_9_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_561 = $signed(hiddenLayers_0_3) * $signed(io_midAndOutputWeights_9_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_562 = $signed(hiddenLayers_0_4) * $signed(io_midAndOutputWeights_9_4); // @[FixedPointTypeClass.scala 43:59]
  assign _T_563 = $signed(hiddenLayers_0_5) * $signed(io_midAndOutputWeights_9_5); // @[FixedPointTypeClass.scala 43:59]
  assign _T_564 = $signed(hiddenLayers_0_6) * $signed(io_midAndOutputWeights_9_6); // @[FixedPointTypeClass.scala 43:59]
  assign _T_565 = $signed(hiddenLayers_0_7) * $signed(io_midAndOutputWeights_9_7); // @[FixedPointTypeClass.scala 43:59]
  assign _T_566 = $signed(hiddenLayers_0_8) * $signed(io_midAndOutputWeights_9_8); // @[FixedPointTypeClass.scala 43:59]
  assign _T_567 = $signed(hiddenLayers_0_9) * $signed(io_midAndOutputWeights_9_9); // @[FixedPointTypeClass.scala 43:59]
  assign _T_569 = $signed(_T_558) + $signed(_T_559); // @[FixedPointTypeClass.scala 21:58]
  assign _T_570 = $signed(_T_569); // @[FixedPointTypeClass.scala 21:58]
  assign _T_572 = $signed(_T_570) + $signed(_T_560); // @[FixedPointTypeClass.scala 21:58]
  assign _T_573 = $signed(_T_572); // @[FixedPointTypeClass.scala 21:58]
  assign _T_575 = $signed(_T_573) + $signed(_T_561); // @[FixedPointTypeClass.scala 21:58]
  assign _T_576 = $signed(_T_575); // @[FixedPointTypeClass.scala 21:58]
  assign _T_578 = $signed(_T_576) + $signed(_T_562); // @[FixedPointTypeClass.scala 21:58]
  assign _T_579 = $signed(_T_578); // @[FixedPointTypeClass.scala 21:58]
  assign _T_581 = $signed(_T_579) + $signed(_T_563); // @[FixedPointTypeClass.scala 21:58]
  assign _T_582 = $signed(_T_581); // @[FixedPointTypeClass.scala 21:58]
  assign _T_584 = $signed(_T_582) + $signed(_T_564); // @[FixedPointTypeClass.scala 21:58]
  assign _T_585 = $signed(_T_584); // @[FixedPointTypeClass.scala 21:58]
  assign _T_587 = $signed(_T_585) + $signed(_T_565); // @[FixedPointTypeClass.scala 21:58]
  assign _T_588 = $signed(_T_587); // @[FixedPointTypeClass.scala 21:58]
  assign _T_590 = $signed(_T_588) + $signed(_T_566); // @[FixedPointTypeClass.scala 21:58]
  assign _T_591 = $signed(_T_590); // @[FixedPointTypeClass.scala 21:58]
  assign _T_593 = $signed(_T_591) + $signed(_T_567); // @[FixedPointTypeClass.scala 21:58]
  assign _T_594 = $signed(_T_593); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_79 = {{8{io_biasVecs_1_9[31]}},io_biasVecs_1_9}; // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_80 = $signed(_GEN_79) << 8; // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_81 = {{24{_GEN_80[39]}},_GEN_80}; // @[FixedPointTypeClass.scala 21:58]
  assign _T_596 = $signed(_T_594) + $signed(_GEN_81); // @[FixedPointTypeClass.scala 21:58]
  assign _T_597 = $signed(_T_596); // @[FixedPointTypeClass.scala 21:58]
  assign _T_598 = $signed(_T_597) > $signed(64'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign _T_599 = _T_598 ? $signed(_T_597) : $signed(64'sh0); // @[neuralNet.scala 59:32]
  assign _GEN_82 = _T_221[63:8]; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  assign _GEN_83 = _GEN_82[31:0]; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  assign hiddenLayers_1_0 = $signed(_GEN_83); // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  assign _T_600 = $signed(hiddenLayers_1_0) * $signed(io_midAndOutputWeights_10_0); // @[FixedPointTypeClass.scala 43:59]
  assign _GEN_84 = _T_263[63:8]; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  assign _GEN_85 = _GEN_84[31:0]; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  assign hiddenLayers_1_1 = $signed(_GEN_85); // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  assign _T_601 = $signed(hiddenLayers_1_1) * $signed(io_midAndOutputWeights_10_1); // @[FixedPointTypeClass.scala 43:59]
  assign _GEN_86 = _T_305[63:8]; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  assign _GEN_87 = _GEN_86[31:0]; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  assign hiddenLayers_1_2 = $signed(_GEN_87); // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  assign _T_602 = $signed(hiddenLayers_1_2) * $signed(io_midAndOutputWeights_10_2); // @[FixedPointTypeClass.scala 43:59]
  assign _GEN_88 = _T_347[63:8]; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  assign _GEN_89 = _GEN_88[31:0]; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  assign hiddenLayers_1_3 = $signed(_GEN_89); // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  assign _T_603 = $signed(hiddenLayers_1_3) * $signed(io_midAndOutputWeights_10_3); // @[FixedPointTypeClass.scala 43:59]
  assign _GEN_90 = _T_389[63:8]; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  assign _GEN_91 = _GEN_90[31:0]; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  assign hiddenLayers_1_4 = $signed(_GEN_91); // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  assign _T_604 = $signed(hiddenLayers_1_4) * $signed(io_midAndOutputWeights_10_4); // @[FixedPointTypeClass.scala 43:59]
  assign _GEN_92 = _T_431[63:8]; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  assign _GEN_93 = _GEN_92[31:0]; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  assign hiddenLayers_1_5 = $signed(_GEN_93); // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  assign _T_605 = $signed(hiddenLayers_1_5) * $signed(io_midAndOutputWeights_10_5); // @[FixedPointTypeClass.scala 43:59]
  assign _GEN_94 = _T_473[63:8]; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  assign _GEN_95 = _GEN_94[31:0]; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  assign hiddenLayers_1_6 = $signed(_GEN_95); // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  assign _T_606 = $signed(hiddenLayers_1_6) * $signed(io_midAndOutputWeights_10_6); // @[FixedPointTypeClass.scala 43:59]
  assign _GEN_96 = _T_515[63:8]; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  assign _GEN_97 = _GEN_96[31:0]; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  assign hiddenLayers_1_7 = $signed(_GEN_97); // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  assign _T_607 = $signed(hiddenLayers_1_7) * $signed(io_midAndOutputWeights_10_7); // @[FixedPointTypeClass.scala 43:59]
  assign _GEN_98 = _T_557[63:8]; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  assign _GEN_99 = _GEN_98[31:0]; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  assign hiddenLayers_1_8 = $signed(_GEN_99); // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  assign _T_608 = $signed(hiddenLayers_1_8) * $signed(io_midAndOutputWeights_10_8); // @[FixedPointTypeClass.scala 43:59]
  assign _GEN_100 = _T_599[63:8]; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  assign _GEN_101 = _GEN_100[31:0]; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  assign hiddenLayers_1_9 = $signed(_GEN_101); // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  assign _T_609 = $signed(hiddenLayers_1_9) * $signed(io_midAndOutputWeights_10_9); // @[FixedPointTypeClass.scala 43:59]
  assign _T_611 = $signed(_T_600) + $signed(_T_601); // @[FixedPointTypeClass.scala 21:58]
  assign _T_612 = $signed(_T_611); // @[FixedPointTypeClass.scala 21:58]
  assign _T_614 = $signed(_T_612) + $signed(_T_602); // @[FixedPointTypeClass.scala 21:58]
  assign _T_615 = $signed(_T_614); // @[FixedPointTypeClass.scala 21:58]
  assign _T_617 = $signed(_T_615) + $signed(_T_603); // @[FixedPointTypeClass.scala 21:58]
  assign _T_618 = $signed(_T_617); // @[FixedPointTypeClass.scala 21:58]
  assign _T_620 = $signed(_T_618) + $signed(_T_604); // @[FixedPointTypeClass.scala 21:58]
  assign _T_621 = $signed(_T_620); // @[FixedPointTypeClass.scala 21:58]
  assign _T_623 = $signed(_T_621) + $signed(_T_605); // @[FixedPointTypeClass.scala 21:58]
  assign _T_624 = $signed(_T_623); // @[FixedPointTypeClass.scala 21:58]
  assign _T_626 = $signed(_T_624) + $signed(_T_606); // @[FixedPointTypeClass.scala 21:58]
  assign _T_627 = $signed(_T_626); // @[FixedPointTypeClass.scala 21:58]
  assign _T_629 = $signed(_T_627) + $signed(_T_607); // @[FixedPointTypeClass.scala 21:58]
  assign _T_630 = $signed(_T_629); // @[FixedPointTypeClass.scala 21:58]
  assign _T_632 = $signed(_T_630) + $signed(_T_608); // @[FixedPointTypeClass.scala 21:58]
  assign _T_633 = $signed(_T_632); // @[FixedPointTypeClass.scala 21:58]
  assign _T_635 = $signed(_T_633) + $signed(_T_609); // @[FixedPointTypeClass.scala 21:58]
  assign _T_636 = $signed(_T_635); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_102 = {{8{io_biasVecs_2_0[31]}},io_biasVecs_2_0}; // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_103 = $signed(_GEN_102) << 8; // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_104 = {{24{_GEN_103[39]}},_GEN_103}; // @[FixedPointTypeClass.scala 21:58]
  assign _T_638 = $signed(_T_636) + $signed(_GEN_104); // @[FixedPointTypeClass.scala 21:58]
  assign _T_639 = $signed(_T_638); // @[FixedPointTypeClass.scala 21:58]
  assign _T_640 = $signed(_T_639) > $signed(64'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign _T_641 = _T_640 ? $signed(_T_639) : $signed(64'sh0); // @[neuralNet.scala 59:32]
  assign _T_642 = $signed(hiddenLayers_1_0) * $signed(io_midAndOutputWeights_11_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_643 = $signed(hiddenLayers_1_1) * $signed(io_midAndOutputWeights_11_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_644 = $signed(hiddenLayers_1_2) * $signed(io_midAndOutputWeights_11_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_645 = $signed(hiddenLayers_1_3) * $signed(io_midAndOutputWeights_11_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_646 = $signed(hiddenLayers_1_4) * $signed(io_midAndOutputWeights_11_4); // @[FixedPointTypeClass.scala 43:59]
  assign _T_647 = $signed(hiddenLayers_1_5) * $signed(io_midAndOutputWeights_11_5); // @[FixedPointTypeClass.scala 43:59]
  assign _T_648 = $signed(hiddenLayers_1_6) * $signed(io_midAndOutputWeights_11_6); // @[FixedPointTypeClass.scala 43:59]
  assign _T_649 = $signed(hiddenLayers_1_7) * $signed(io_midAndOutputWeights_11_7); // @[FixedPointTypeClass.scala 43:59]
  assign _T_650 = $signed(hiddenLayers_1_8) * $signed(io_midAndOutputWeights_11_8); // @[FixedPointTypeClass.scala 43:59]
  assign _T_651 = $signed(hiddenLayers_1_9) * $signed(io_midAndOutputWeights_11_9); // @[FixedPointTypeClass.scala 43:59]
  assign _T_653 = $signed(_T_642) + $signed(_T_643); // @[FixedPointTypeClass.scala 21:58]
  assign _T_654 = $signed(_T_653); // @[FixedPointTypeClass.scala 21:58]
  assign _T_656 = $signed(_T_654) + $signed(_T_644); // @[FixedPointTypeClass.scala 21:58]
  assign _T_657 = $signed(_T_656); // @[FixedPointTypeClass.scala 21:58]
  assign _T_659 = $signed(_T_657) + $signed(_T_645); // @[FixedPointTypeClass.scala 21:58]
  assign _T_660 = $signed(_T_659); // @[FixedPointTypeClass.scala 21:58]
  assign _T_662 = $signed(_T_660) + $signed(_T_646); // @[FixedPointTypeClass.scala 21:58]
  assign _T_663 = $signed(_T_662); // @[FixedPointTypeClass.scala 21:58]
  assign _T_665 = $signed(_T_663) + $signed(_T_647); // @[FixedPointTypeClass.scala 21:58]
  assign _T_666 = $signed(_T_665); // @[FixedPointTypeClass.scala 21:58]
  assign _T_668 = $signed(_T_666) + $signed(_T_648); // @[FixedPointTypeClass.scala 21:58]
  assign _T_669 = $signed(_T_668); // @[FixedPointTypeClass.scala 21:58]
  assign _T_671 = $signed(_T_669) + $signed(_T_649); // @[FixedPointTypeClass.scala 21:58]
  assign _T_672 = $signed(_T_671); // @[FixedPointTypeClass.scala 21:58]
  assign _T_674 = $signed(_T_672) + $signed(_T_650); // @[FixedPointTypeClass.scala 21:58]
  assign _T_675 = $signed(_T_674); // @[FixedPointTypeClass.scala 21:58]
  assign _T_677 = $signed(_T_675) + $signed(_T_651); // @[FixedPointTypeClass.scala 21:58]
  assign _T_678 = $signed(_T_677); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_105 = {{8{io_biasVecs_2_1[31]}},io_biasVecs_2_1}; // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_106 = $signed(_GEN_105) << 8; // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_107 = {{24{_GEN_106[39]}},_GEN_106}; // @[FixedPointTypeClass.scala 21:58]
  assign _T_680 = $signed(_T_678) + $signed(_GEN_107); // @[FixedPointTypeClass.scala 21:58]
  assign _T_681 = $signed(_T_680); // @[FixedPointTypeClass.scala 21:58]
  assign _T_682 = $signed(_T_681) > $signed(64'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign _T_683 = _T_682 ? $signed(_T_681) : $signed(64'sh0); // @[neuralNet.scala 59:32]
  assign _T_684 = $signed(hiddenLayers_1_0) * $signed(io_midAndOutputWeights_12_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_685 = $signed(hiddenLayers_1_1) * $signed(io_midAndOutputWeights_12_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_686 = $signed(hiddenLayers_1_2) * $signed(io_midAndOutputWeights_12_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_687 = $signed(hiddenLayers_1_3) * $signed(io_midAndOutputWeights_12_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_688 = $signed(hiddenLayers_1_4) * $signed(io_midAndOutputWeights_12_4); // @[FixedPointTypeClass.scala 43:59]
  assign _T_689 = $signed(hiddenLayers_1_5) * $signed(io_midAndOutputWeights_12_5); // @[FixedPointTypeClass.scala 43:59]
  assign _T_690 = $signed(hiddenLayers_1_6) * $signed(io_midAndOutputWeights_12_6); // @[FixedPointTypeClass.scala 43:59]
  assign _T_691 = $signed(hiddenLayers_1_7) * $signed(io_midAndOutputWeights_12_7); // @[FixedPointTypeClass.scala 43:59]
  assign _T_692 = $signed(hiddenLayers_1_8) * $signed(io_midAndOutputWeights_12_8); // @[FixedPointTypeClass.scala 43:59]
  assign _T_693 = $signed(hiddenLayers_1_9) * $signed(io_midAndOutputWeights_12_9); // @[FixedPointTypeClass.scala 43:59]
  assign _T_695 = $signed(_T_684) + $signed(_T_685); // @[FixedPointTypeClass.scala 21:58]
  assign _T_696 = $signed(_T_695); // @[FixedPointTypeClass.scala 21:58]
  assign _T_698 = $signed(_T_696) + $signed(_T_686); // @[FixedPointTypeClass.scala 21:58]
  assign _T_699 = $signed(_T_698); // @[FixedPointTypeClass.scala 21:58]
  assign _T_701 = $signed(_T_699) + $signed(_T_687); // @[FixedPointTypeClass.scala 21:58]
  assign _T_702 = $signed(_T_701); // @[FixedPointTypeClass.scala 21:58]
  assign _T_704 = $signed(_T_702) + $signed(_T_688); // @[FixedPointTypeClass.scala 21:58]
  assign _T_705 = $signed(_T_704); // @[FixedPointTypeClass.scala 21:58]
  assign _T_707 = $signed(_T_705) + $signed(_T_689); // @[FixedPointTypeClass.scala 21:58]
  assign _T_708 = $signed(_T_707); // @[FixedPointTypeClass.scala 21:58]
  assign _T_710 = $signed(_T_708) + $signed(_T_690); // @[FixedPointTypeClass.scala 21:58]
  assign _T_711 = $signed(_T_710); // @[FixedPointTypeClass.scala 21:58]
  assign _T_713 = $signed(_T_711) + $signed(_T_691); // @[FixedPointTypeClass.scala 21:58]
  assign _T_714 = $signed(_T_713); // @[FixedPointTypeClass.scala 21:58]
  assign _T_716 = $signed(_T_714) + $signed(_T_692); // @[FixedPointTypeClass.scala 21:58]
  assign _T_717 = $signed(_T_716); // @[FixedPointTypeClass.scala 21:58]
  assign _T_719 = $signed(_T_717) + $signed(_T_693); // @[FixedPointTypeClass.scala 21:58]
  assign _T_720 = $signed(_T_719); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_108 = {{8{io_biasVecs_2_2[31]}},io_biasVecs_2_2}; // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_109 = $signed(_GEN_108) << 8; // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_110 = {{24{_GEN_109[39]}},_GEN_109}; // @[FixedPointTypeClass.scala 21:58]
  assign _T_722 = $signed(_T_720) + $signed(_GEN_110); // @[FixedPointTypeClass.scala 21:58]
  assign _T_723 = $signed(_T_722); // @[FixedPointTypeClass.scala 21:58]
  assign _T_724 = $signed(_T_723) > $signed(64'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign _T_725 = _T_724 ? $signed(_T_723) : $signed(64'sh0); // @[neuralNet.scala 59:32]
  assign _T_726 = $signed(hiddenLayers_1_0) * $signed(io_midAndOutputWeights_13_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_727 = $signed(hiddenLayers_1_1) * $signed(io_midAndOutputWeights_13_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_728 = $signed(hiddenLayers_1_2) * $signed(io_midAndOutputWeights_13_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_729 = $signed(hiddenLayers_1_3) * $signed(io_midAndOutputWeights_13_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_730 = $signed(hiddenLayers_1_4) * $signed(io_midAndOutputWeights_13_4); // @[FixedPointTypeClass.scala 43:59]
  assign _T_731 = $signed(hiddenLayers_1_5) * $signed(io_midAndOutputWeights_13_5); // @[FixedPointTypeClass.scala 43:59]
  assign _T_732 = $signed(hiddenLayers_1_6) * $signed(io_midAndOutputWeights_13_6); // @[FixedPointTypeClass.scala 43:59]
  assign _T_733 = $signed(hiddenLayers_1_7) * $signed(io_midAndOutputWeights_13_7); // @[FixedPointTypeClass.scala 43:59]
  assign _T_734 = $signed(hiddenLayers_1_8) * $signed(io_midAndOutputWeights_13_8); // @[FixedPointTypeClass.scala 43:59]
  assign _T_735 = $signed(hiddenLayers_1_9) * $signed(io_midAndOutputWeights_13_9); // @[FixedPointTypeClass.scala 43:59]
  assign _T_737 = $signed(_T_726) + $signed(_T_727); // @[FixedPointTypeClass.scala 21:58]
  assign _T_738 = $signed(_T_737); // @[FixedPointTypeClass.scala 21:58]
  assign _T_740 = $signed(_T_738) + $signed(_T_728); // @[FixedPointTypeClass.scala 21:58]
  assign _T_741 = $signed(_T_740); // @[FixedPointTypeClass.scala 21:58]
  assign _T_743 = $signed(_T_741) + $signed(_T_729); // @[FixedPointTypeClass.scala 21:58]
  assign _T_744 = $signed(_T_743); // @[FixedPointTypeClass.scala 21:58]
  assign _T_746 = $signed(_T_744) + $signed(_T_730); // @[FixedPointTypeClass.scala 21:58]
  assign _T_747 = $signed(_T_746); // @[FixedPointTypeClass.scala 21:58]
  assign _T_749 = $signed(_T_747) + $signed(_T_731); // @[FixedPointTypeClass.scala 21:58]
  assign _T_750 = $signed(_T_749); // @[FixedPointTypeClass.scala 21:58]
  assign _T_752 = $signed(_T_750) + $signed(_T_732); // @[FixedPointTypeClass.scala 21:58]
  assign _T_753 = $signed(_T_752); // @[FixedPointTypeClass.scala 21:58]
  assign _T_755 = $signed(_T_753) + $signed(_T_733); // @[FixedPointTypeClass.scala 21:58]
  assign _T_756 = $signed(_T_755); // @[FixedPointTypeClass.scala 21:58]
  assign _T_758 = $signed(_T_756) + $signed(_T_734); // @[FixedPointTypeClass.scala 21:58]
  assign _T_759 = $signed(_T_758); // @[FixedPointTypeClass.scala 21:58]
  assign _T_761 = $signed(_T_759) + $signed(_T_735); // @[FixedPointTypeClass.scala 21:58]
  assign _T_762 = $signed(_T_761); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_111 = {{8{io_biasVecs_2_3[31]}},io_biasVecs_2_3}; // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_112 = $signed(_GEN_111) << 8; // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_113 = {{24{_GEN_112[39]}},_GEN_112}; // @[FixedPointTypeClass.scala 21:58]
  assign _T_764 = $signed(_T_762) + $signed(_GEN_113); // @[FixedPointTypeClass.scala 21:58]
  assign _T_765 = $signed(_T_764); // @[FixedPointTypeClass.scala 21:58]
  assign _T_766 = $signed(_T_765) > $signed(64'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign _T_767 = _T_766 ? $signed(_T_765) : $signed(64'sh0); // @[neuralNet.scala 59:32]
  assign _T_768 = $signed(hiddenLayers_1_0) * $signed(io_midAndOutputWeights_14_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_769 = $signed(hiddenLayers_1_1) * $signed(io_midAndOutputWeights_14_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_770 = $signed(hiddenLayers_1_2) * $signed(io_midAndOutputWeights_14_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_771 = $signed(hiddenLayers_1_3) * $signed(io_midAndOutputWeights_14_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_772 = $signed(hiddenLayers_1_4) * $signed(io_midAndOutputWeights_14_4); // @[FixedPointTypeClass.scala 43:59]
  assign _T_773 = $signed(hiddenLayers_1_5) * $signed(io_midAndOutputWeights_14_5); // @[FixedPointTypeClass.scala 43:59]
  assign _T_774 = $signed(hiddenLayers_1_6) * $signed(io_midAndOutputWeights_14_6); // @[FixedPointTypeClass.scala 43:59]
  assign _T_775 = $signed(hiddenLayers_1_7) * $signed(io_midAndOutputWeights_14_7); // @[FixedPointTypeClass.scala 43:59]
  assign _T_776 = $signed(hiddenLayers_1_8) * $signed(io_midAndOutputWeights_14_8); // @[FixedPointTypeClass.scala 43:59]
  assign _T_777 = $signed(hiddenLayers_1_9) * $signed(io_midAndOutputWeights_14_9); // @[FixedPointTypeClass.scala 43:59]
  assign _T_779 = $signed(_T_768) + $signed(_T_769); // @[FixedPointTypeClass.scala 21:58]
  assign _T_780 = $signed(_T_779); // @[FixedPointTypeClass.scala 21:58]
  assign _T_782 = $signed(_T_780) + $signed(_T_770); // @[FixedPointTypeClass.scala 21:58]
  assign _T_783 = $signed(_T_782); // @[FixedPointTypeClass.scala 21:58]
  assign _T_785 = $signed(_T_783) + $signed(_T_771); // @[FixedPointTypeClass.scala 21:58]
  assign _T_786 = $signed(_T_785); // @[FixedPointTypeClass.scala 21:58]
  assign _T_788 = $signed(_T_786) + $signed(_T_772); // @[FixedPointTypeClass.scala 21:58]
  assign _T_789 = $signed(_T_788); // @[FixedPointTypeClass.scala 21:58]
  assign _T_791 = $signed(_T_789) + $signed(_T_773); // @[FixedPointTypeClass.scala 21:58]
  assign _T_792 = $signed(_T_791); // @[FixedPointTypeClass.scala 21:58]
  assign _T_794 = $signed(_T_792) + $signed(_T_774); // @[FixedPointTypeClass.scala 21:58]
  assign _T_795 = $signed(_T_794); // @[FixedPointTypeClass.scala 21:58]
  assign _T_797 = $signed(_T_795) + $signed(_T_775); // @[FixedPointTypeClass.scala 21:58]
  assign _T_798 = $signed(_T_797); // @[FixedPointTypeClass.scala 21:58]
  assign _T_800 = $signed(_T_798) + $signed(_T_776); // @[FixedPointTypeClass.scala 21:58]
  assign _T_801 = $signed(_T_800); // @[FixedPointTypeClass.scala 21:58]
  assign _T_803 = $signed(_T_801) + $signed(_T_777); // @[FixedPointTypeClass.scala 21:58]
  assign _T_804 = $signed(_T_803); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_114 = {{8{io_biasVecs_2_4[31]}},io_biasVecs_2_4}; // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_115 = $signed(_GEN_114) << 8; // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_116 = {{24{_GEN_115[39]}},_GEN_115}; // @[FixedPointTypeClass.scala 21:58]
  assign _T_806 = $signed(_T_804) + $signed(_GEN_116); // @[FixedPointTypeClass.scala 21:58]
  assign _T_807 = $signed(_T_806); // @[FixedPointTypeClass.scala 21:58]
  assign _T_808 = $signed(_T_807) > $signed(64'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign _T_809 = _T_808 ? $signed(_T_807) : $signed(64'sh0); // @[neuralNet.scala 59:32]
  assign _T_810 = $signed(hiddenLayers_1_0) * $signed(io_midAndOutputWeights_15_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_811 = $signed(hiddenLayers_1_1) * $signed(io_midAndOutputWeights_15_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_812 = $signed(hiddenLayers_1_2) * $signed(io_midAndOutputWeights_15_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_813 = $signed(hiddenLayers_1_3) * $signed(io_midAndOutputWeights_15_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_814 = $signed(hiddenLayers_1_4) * $signed(io_midAndOutputWeights_15_4); // @[FixedPointTypeClass.scala 43:59]
  assign _T_815 = $signed(hiddenLayers_1_5) * $signed(io_midAndOutputWeights_15_5); // @[FixedPointTypeClass.scala 43:59]
  assign _T_816 = $signed(hiddenLayers_1_6) * $signed(io_midAndOutputWeights_15_6); // @[FixedPointTypeClass.scala 43:59]
  assign _T_817 = $signed(hiddenLayers_1_7) * $signed(io_midAndOutputWeights_15_7); // @[FixedPointTypeClass.scala 43:59]
  assign _T_818 = $signed(hiddenLayers_1_8) * $signed(io_midAndOutputWeights_15_8); // @[FixedPointTypeClass.scala 43:59]
  assign _T_819 = $signed(hiddenLayers_1_9) * $signed(io_midAndOutputWeights_15_9); // @[FixedPointTypeClass.scala 43:59]
  assign _T_821 = $signed(_T_810) + $signed(_T_811); // @[FixedPointTypeClass.scala 21:58]
  assign _T_822 = $signed(_T_821); // @[FixedPointTypeClass.scala 21:58]
  assign _T_824 = $signed(_T_822) + $signed(_T_812); // @[FixedPointTypeClass.scala 21:58]
  assign _T_825 = $signed(_T_824); // @[FixedPointTypeClass.scala 21:58]
  assign _T_827 = $signed(_T_825) + $signed(_T_813); // @[FixedPointTypeClass.scala 21:58]
  assign _T_828 = $signed(_T_827); // @[FixedPointTypeClass.scala 21:58]
  assign _T_830 = $signed(_T_828) + $signed(_T_814); // @[FixedPointTypeClass.scala 21:58]
  assign _T_831 = $signed(_T_830); // @[FixedPointTypeClass.scala 21:58]
  assign _T_833 = $signed(_T_831) + $signed(_T_815); // @[FixedPointTypeClass.scala 21:58]
  assign _T_834 = $signed(_T_833); // @[FixedPointTypeClass.scala 21:58]
  assign _T_836 = $signed(_T_834) + $signed(_T_816); // @[FixedPointTypeClass.scala 21:58]
  assign _T_837 = $signed(_T_836); // @[FixedPointTypeClass.scala 21:58]
  assign _T_839 = $signed(_T_837) + $signed(_T_817); // @[FixedPointTypeClass.scala 21:58]
  assign _T_840 = $signed(_T_839); // @[FixedPointTypeClass.scala 21:58]
  assign _T_842 = $signed(_T_840) + $signed(_T_818); // @[FixedPointTypeClass.scala 21:58]
  assign _T_843 = $signed(_T_842); // @[FixedPointTypeClass.scala 21:58]
  assign _T_845 = $signed(_T_843) + $signed(_T_819); // @[FixedPointTypeClass.scala 21:58]
  assign _T_846 = $signed(_T_845); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_117 = {{8{io_biasVecs_2_5[31]}},io_biasVecs_2_5}; // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_118 = $signed(_GEN_117) << 8; // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_119 = {{24{_GEN_118[39]}},_GEN_118}; // @[FixedPointTypeClass.scala 21:58]
  assign _T_848 = $signed(_T_846) + $signed(_GEN_119); // @[FixedPointTypeClass.scala 21:58]
  assign _T_849 = $signed(_T_848); // @[FixedPointTypeClass.scala 21:58]
  assign _T_850 = $signed(_T_849) > $signed(64'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign _T_851 = _T_850 ? $signed(_T_849) : $signed(64'sh0); // @[neuralNet.scala 59:32]
  assign _T_852 = $signed(hiddenLayers_1_0) * $signed(io_midAndOutputWeights_16_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_853 = $signed(hiddenLayers_1_1) * $signed(io_midAndOutputWeights_16_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_854 = $signed(hiddenLayers_1_2) * $signed(io_midAndOutputWeights_16_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_855 = $signed(hiddenLayers_1_3) * $signed(io_midAndOutputWeights_16_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_856 = $signed(hiddenLayers_1_4) * $signed(io_midAndOutputWeights_16_4); // @[FixedPointTypeClass.scala 43:59]
  assign _T_857 = $signed(hiddenLayers_1_5) * $signed(io_midAndOutputWeights_16_5); // @[FixedPointTypeClass.scala 43:59]
  assign _T_858 = $signed(hiddenLayers_1_6) * $signed(io_midAndOutputWeights_16_6); // @[FixedPointTypeClass.scala 43:59]
  assign _T_859 = $signed(hiddenLayers_1_7) * $signed(io_midAndOutputWeights_16_7); // @[FixedPointTypeClass.scala 43:59]
  assign _T_860 = $signed(hiddenLayers_1_8) * $signed(io_midAndOutputWeights_16_8); // @[FixedPointTypeClass.scala 43:59]
  assign _T_861 = $signed(hiddenLayers_1_9) * $signed(io_midAndOutputWeights_16_9); // @[FixedPointTypeClass.scala 43:59]
  assign _T_863 = $signed(_T_852) + $signed(_T_853); // @[FixedPointTypeClass.scala 21:58]
  assign _T_864 = $signed(_T_863); // @[FixedPointTypeClass.scala 21:58]
  assign _T_866 = $signed(_T_864) + $signed(_T_854); // @[FixedPointTypeClass.scala 21:58]
  assign _T_867 = $signed(_T_866); // @[FixedPointTypeClass.scala 21:58]
  assign _T_869 = $signed(_T_867) + $signed(_T_855); // @[FixedPointTypeClass.scala 21:58]
  assign _T_870 = $signed(_T_869); // @[FixedPointTypeClass.scala 21:58]
  assign _T_872 = $signed(_T_870) + $signed(_T_856); // @[FixedPointTypeClass.scala 21:58]
  assign _T_873 = $signed(_T_872); // @[FixedPointTypeClass.scala 21:58]
  assign _T_875 = $signed(_T_873) + $signed(_T_857); // @[FixedPointTypeClass.scala 21:58]
  assign _T_876 = $signed(_T_875); // @[FixedPointTypeClass.scala 21:58]
  assign _T_878 = $signed(_T_876) + $signed(_T_858); // @[FixedPointTypeClass.scala 21:58]
  assign _T_879 = $signed(_T_878); // @[FixedPointTypeClass.scala 21:58]
  assign _T_881 = $signed(_T_879) + $signed(_T_859); // @[FixedPointTypeClass.scala 21:58]
  assign _T_882 = $signed(_T_881); // @[FixedPointTypeClass.scala 21:58]
  assign _T_884 = $signed(_T_882) + $signed(_T_860); // @[FixedPointTypeClass.scala 21:58]
  assign _T_885 = $signed(_T_884); // @[FixedPointTypeClass.scala 21:58]
  assign _T_887 = $signed(_T_885) + $signed(_T_861); // @[FixedPointTypeClass.scala 21:58]
  assign _T_888 = $signed(_T_887); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_120 = {{8{io_biasVecs_2_6[31]}},io_biasVecs_2_6}; // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_121 = $signed(_GEN_120) << 8; // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_122 = {{24{_GEN_121[39]}},_GEN_121}; // @[FixedPointTypeClass.scala 21:58]
  assign _T_890 = $signed(_T_888) + $signed(_GEN_122); // @[FixedPointTypeClass.scala 21:58]
  assign _T_891 = $signed(_T_890); // @[FixedPointTypeClass.scala 21:58]
  assign _T_892 = $signed(_T_891) > $signed(64'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign _T_893 = _T_892 ? $signed(_T_891) : $signed(64'sh0); // @[neuralNet.scala 59:32]
  assign _T_894 = $signed(hiddenLayers_1_0) * $signed(io_midAndOutputWeights_17_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_895 = $signed(hiddenLayers_1_1) * $signed(io_midAndOutputWeights_17_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_896 = $signed(hiddenLayers_1_2) * $signed(io_midAndOutputWeights_17_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_897 = $signed(hiddenLayers_1_3) * $signed(io_midAndOutputWeights_17_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_898 = $signed(hiddenLayers_1_4) * $signed(io_midAndOutputWeights_17_4); // @[FixedPointTypeClass.scala 43:59]
  assign _T_899 = $signed(hiddenLayers_1_5) * $signed(io_midAndOutputWeights_17_5); // @[FixedPointTypeClass.scala 43:59]
  assign _T_900 = $signed(hiddenLayers_1_6) * $signed(io_midAndOutputWeights_17_6); // @[FixedPointTypeClass.scala 43:59]
  assign _T_901 = $signed(hiddenLayers_1_7) * $signed(io_midAndOutputWeights_17_7); // @[FixedPointTypeClass.scala 43:59]
  assign _T_902 = $signed(hiddenLayers_1_8) * $signed(io_midAndOutputWeights_17_8); // @[FixedPointTypeClass.scala 43:59]
  assign _T_903 = $signed(hiddenLayers_1_9) * $signed(io_midAndOutputWeights_17_9); // @[FixedPointTypeClass.scala 43:59]
  assign _T_905 = $signed(_T_894) + $signed(_T_895); // @[FixedPointTypeClass.scala 21:58]
  assign _T_906 = $signed(_T_905); // @[FixedPointTypeClass.scala 21:58]
  assign _T_908 = $signed(_T_906) + $signed(_T_896); // @[FixedPointTypeClass.scala 21:58]
  assign _T_909 = $signed(_T_908); // @[FixedPointTypeClass.scala 21:58]
  assign _T_911 = $signed(_T_909) + $signed(_T_897); // @[FixedPointTypeClass.scala 21:58]
  assign _T_912 = $signed(_T_911); // @[FixedPointTypeClass.scala 21:58]
  assign _T_914 = $signed(_T_912) + $signed(_T_898); // @[FixedPointTypeClass.scala 21:58]
  assign _T_915 = $signed(_T_914); // @[FixedPointTypeClass.scala 21:58]
  assign _T_917 = $signed(_T_915) + $signed(_T_899); // @[FixedPointTypeClass.scala 21:58]
  assign _T_918 = $signed(_T_917); // @[FixedPointTypeClass.scala 21:58]
  assign _T_920 = $signed(_T_918) + $signed(_T_900); // @[FixedPointTypeClass.scala 21:58]
  assign _T_921 = $signed(_T_920); // @[FixedPointTypeClass.scala 21:58]
  assign _T_923 = $signed(_T_921) + $signed(_T_901); // @[FixedPointTypeClass.scala 21:58]
  assign _T_924 = $signed(_T_923); // @[FixedPointTypeClass.scala 21:58]
  assign _T_926 = $signed(_T_924) + $signed(_T_902); // @[FixedPointTypeClass.scala 21:58]
  assign _T_927 = $signed(_T_926); // @[FixedPointTypeClass.scala 21:58]
  assign _T_929 = $signed(_T_927) + $signed(_T_903); // @[FixedPointTypeClass.scala 21:58]
  assign _T_930 = $signed(_T_929); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_123 = {{8{io_biasVecs_2_7[31]}},io_biasVecs_2_7}; // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_124 = $signed(_GEN_123) << 8; // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_125 = {{24{_GEN_124[39]}},_GEN_124}; // @[FixedPointTypeClass.scala 21:58]
  assign _T_932 = $signed(_T_930) + $signed(_GEN_125); // @[FixedPointTypeClass.scala 21:58]
  assign _T_933 = $signed(_T_932); // @[FixedPointTypeClass.scala 21:58]
  assign _T_934 = $signed(_T_933) > $signed(64'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign _T_935 = _T_934 ? $signed(_T_933) : $signed(64'sh0); // @[neuralNet.scala 59:32]
  assign _T_936 = $signed(hiddenLayers_1_0) * $signed(io_midAndOutputWeights_18_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_937 = $signed(hiddenLayers_1_1) * $signed(io_midAndOutputWeights_18_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_938 = $signed(hiddenLayers_1_2) * $signed(io_midAndOutputWeights_18_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_939 = $signed(hiddenLayers_1_3) * $signed(io_midAndOutputWeights_18_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_940 = $signed(hiddenLayers_1_4) * $signed(io_midAndOutputWeights_18_4); // @[FixedPointTypeClass.scala 43:59]
  assign _T_941 = $signed(hiddenLayers_1_5) * $signed(io_midAndOutputWeights_18_5); // @[FixedPointTypeClass.scala 43:59]
  assign _T_942 = $signed(hiddenLayers_1_6) * $signed(io_midAndOutputWeights_18_6); // @[FixedPointTypeClass.scala 43:59]
  assign _T_943 = $signed(hiddenLayers_1_7) * $signed(io_midAndOutputWeights_18_7); // @[FixedPointTypeClass.scala 43:59]
  assign _T_944 = $signed(hiddenLayers_1_8) * $signed(io_midAndOutputWeights_18_8); // @[FixedPointTypeClass.scala 43:59]
  assign _T_945 = $signed(hiddenLayers_1_9) * $signed(io_midAndOutputWeights_18_9); // @[FixedPointTypeClass.scala 43:59]
  assign _T_947 = $signed(_T_936) + $signed(_T_937); // @[FixedPointTypeClass.scala 21:58]
  assign _T_948 = $signed(_T_947); // @[FixedPointTypeClass.scala 21:58]
  assign _T_950 = $signed(_T_948) + $signed(_T_938); // @[FixedPointTypeClass.scala 21:58]
  assign _T_951 = $signed(_T_950); // @[FixedPointTypeClass.scala 21:58]
  assign _T_953 = $signed(_T_951) + $signed(_T_939); // @[FixedPointTypeClass.scala 21:58]
  assign _T_954 = $signed(_T_953); // @[FixedPointTypeClass.scala 21:58]
  assign _T_956 = $signed(_T_954) + $signed(_T_940); // @[FixedPointTypeClass.scala 21:58]
  assign _T_957 = $signed(_T_956); // @[FixedPointTypeClass.scala 21:58]
  assign _T_959 = $signed(_T_957) + $signed(_T_941); // @[FixedPointTypeClass.scala 21:58]
  assign _T_960 = $signed(_T_959); // @[FixedPointTypeClass.scala 21:58]
  assign _T_962 = $signed(_T_960) + $signed(_T_942); // @[FixedPointTypeClass.scala 21:58]
  assign _T_963 = $signed(_T_962); // @[FixedPointTypeClass.scala 21:58]
  assign _T_965 = $signed(_T_963) + $signed(_T_943); // @[FixedPointTypeClass.scala 21:58]
  assign _T_966 = $signed(_T_965); // @[FixedPointTypeClass.scala 21:58]
  assign _T_968 = $signed(_T_966) + $signed(_T_944); // @[FixedPointTypeClass.scala 21:58]
  assign _T_969 = $signed(_T_968); // @[FixedPointTypeClass.scala 21:58]
  assign _T_971 = $signed(_T_969) + $signed(_T_945); // @[FixedPointTypeClass.scala 21:58]
  assign _T_972 = $signed(_T_971); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_126 = {{8{io_biasVecs_2_8[31]}},io_biasVecs_2_8}; // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_127 = $signed(_GEN_126) << 8; // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_128 = {{24{_GEN_127[39]}},_GEN_127}; // @[FixedPointTypeClass.scala 21:58]
  assign _T_974 = $signed(_T_972) + $signed(_GEN_128); // @[FixedPointTypeClass.scala 21:58]
  assign _T_975 = $signed(_T_974); // @[FixedPointTypeClass.scala 21:58]
  assign _T_976 = $signed(_T_975) > $signed(64'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign _T_977 = _T_976 ? $signed(_T_975) : $signed(64'sh0); // @[neuralNet.scala 59:32]
  assign _T_978 = $signed(hiddenLayers_1_0) * $signed(io_midAndOutputWeights_19_0); // @[FixedPointTypeClass.scala 43:59]
  assign _T_979 = $signed(hiddenLayers_1_1) * $signed(io_midAndOutputWeights_19_1); // @[FixedPointTypeClass.scala 43:59]
  assign _T_980 = $signed(hiddenLayers_1_2) * $signed(io_midAndOutputWeights_19_2); // @[FixedPointTypeClass.scala 43:59]
  assign _T_981 = $signed(hiddenLayers_1_3) * $signed(io_midAndOutputWeights_19_3); // @[FixedPointTypeClass.scala 43:59]
  assign _T_982 = $signed(hiddenLayers_1_4) * $signed(io_midAndOutputWeights_19_4); // @[FixedPointTypeClass.scala 43:59]
  assign _T_983 = $signed(hiddenLayers_1_5) * $signed(io_midAndOutputWeights_19_5); // @[FixedPointTypeClass.scala 43:59]
  assign _T_984 = $signed(hiddenLayers_1_6) * $signed(io_midAndOutputWeights_19_6); // @[FixedPointTypeClass.scala 43:59]
  assign _T_985 = $signed(hiddenLayers_1_7) * $signed(io_midAndOutputWeights_19_7); // @[FixedPointTypeClass.scala 43:59]
  assign _T_986 = $signed(hiddenLayers_1_8) * $signed(io_midAndOutputWeights_19_8); // @[FixedPointTypeClass.scala 43:59]
  assign _T_987 = $signed(hiddenLayers_1_9) * $signed(io_midAndOutputWeights_19_9); // @[FixedPointTypeClass.scala 43:59]
  assign _T_989 = $signed(_T_978) + $signed(_T_979); // @[FixedPointTypeClass.scala 21:58]
  assign _T_990 = $signed(_T_989); // @[FixedPointTypeClass.scala 21:58]
  assign _T_992 = $signed(_T_990) + $signed(_T_980); // @[FixedPointTypeClass.scala 21:58]
  assign _T_993 = $signed(_T_992); // @[FixedPointTypeClass.scala 21:58]
  assign _T_995 = $signed(_T_993) + $signed(_T_981); // @[FixedPointTypeClass.scala 21:58]
  assign _T_996 = $signed(_T_995); // @[FixedPointTypeClass.scala 21:58]
  assign _T_998 = $signed(_T_996) + $signed(_T_982); // @[FixedPointTypeClass.scala 21:58]
  assign _T_999 = $signed(_T_998); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1001 = $signed(_T_999) + $signed(_T_983); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1002 = $signed(_T_1001); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1004 = $signed(_T_1002) + $signed(_T_984); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1005 = $signed(_T_1004); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1007 = $signed(_T_1005) + $signed(_T_985); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1008 = $signed(_T_1007); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1010 = $signed(_T_1008) + $signed(_T_986); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1011 = $signed(_T_1010); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1013 = $signed(_T_1011) + $signed(_T_987); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1014 = $signed(_T_1013); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_129 = {{8{io_biasVecs_2_9[31]}},io_biasVecs_2_9}; // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_130 = $signed(_GEN_129) << 8; // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_131 = {{24{_GEN_130[39]}},_GEN_130}; // @[FixedPointTypeClass.scala 21:58]
  assign _T_1016 = $signed(_T_1014) + $signed(_GEN_131); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1017 = $signed(_T_1016); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1018 = $signed(_T_1017) > $signed(64'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign _T_1019 = _T_1018 ? $signed(_T_1017) : $signed(64'sh0); // @[neuralNet.scala 59:32]
  assign _GEN_132 = _T_641[63:8]; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  assign _GEN_133 = _GEN_132[31:0]; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  assign hiddenLayers_2_0 = $signed(_GEN_133); // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  assign _T_1020 = $signed(hiddenLayers_2_0) * $signed(io_midAndOutputWeights_20_0); // @[FixedPointTypeClass.scala 43:59]
  assign _GEN_134 = _T_683[63:8]; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  assign _GEN_135 = _GEN_134[31:0]; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  assign hiddenLayers_2_1 = $signed(_GEN_135); // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  assign _T_1021 = $signed(hiddenLayers_2_1) * $signed(io_midAndOutputWeights_20_1); // @[FixedPointTypeClass.scala 43:59]
  assign _GEN_136 = _T_725[63:8]; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  assign _GEN_137 = _GEN_136[31:0]; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  assign hiddenLayers_2_2 = $signed(_GEN_137); // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  assign _T_1022 = $signed(hiddenLayers_2_2) * $signed(io_midAndOutputWeights_20_2); // @[FixedPointTypeClass.scala 43:59]
  assign _GEN_138 = _T_767[63:8]; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  assign _GEN_139 = _GEN_138[31:0]; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  assign hiddenLayers_2_3 = $signed(_GEN_139); // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  assign _T_1023 = $signed(hiddenLayers_2_3) * $signed(io_midAndOutputWeights_20_3); // @[FixedPointTypeClass.scala 43:59]
  assign _GEN_140 = _T_809[63:8]; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  assign _GEN_141 = _GEN_140[31:0]; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  assign hiddenLayers_2_4 = $signed(_GEN_141); // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  assign _T_1024 = $signed(hiddenLayers_2_4) * $signed(io_midAndOutputWeights_20_4); // @[FixedPointTypeClass.scala 43:59]
  assign _GEN_142 = _T_851[63:8]; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  assign _GEN_143 = _GEN_142[31:0]; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  assign hiddenLayers_2_5 = $signed(_GEN_143); // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  assign _T_1025 = $signed(hiddenLayers_2_5) * $signed(io_midAndOutputWeights_20_5); // @[FixedPointTypeClass.scala 43:59]
  assign _GEN_144 = _T_893[63:8]; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  assign _GEN_145 = _GEN_144[31:0]; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  assign hiddenLayers_2_6 = $signed(_GEN_145); // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  assign _T_1026 = $signed(hiddenLayers_2_6) * $signed(io_midAndOutputWeights_20_6); // @[FixedPointTypeClass.scala 43:59]
  assign _GEN_146 = _T_935[63:8]; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  assign _GEN_147 = _GEN_146[31:0]; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  assign hiddenLayers_2_7 = $signed(_GEN_147); // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  assign _T_1027 = $signed(hiddenLayers_2_7) * $signed(io_midAndOutputWeights_20_7); // @[FixedPointTypeClass.scala 43:59]
  assign _GEN_148 = _T_977[63:8]; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  assign _GEN_149 = _GEN_148[31:0]; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  assign hiddenLayers_2_8 = $signed(_GEN_149); // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  assign _T_1028 = $signed(hiddenLayers_2_8) * $signed(io_midAndOutputWeights_20_8); // @[FixedPointTypeClass.scala 43:59]
  assign _GEN_150 = _T_1019[63:8]; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  assign _GEN_151 = _GEN_150[31:0]; // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  assign hiddenLayers_2_9 = $signed(_GEN_151); // @[neuralNet.scala 43:26 neuralNet.scala 59:26]
  assign _T_1029 = $signed(hiddenLayers_2_9) * $signed(io_midAndOutputWeights_20_9); // @[FixedPointTypeClass.scala 43:59]
  assign _T_1031 = $signed(_T_1020) + $signed(_T_1021); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1032 = $signed(_T_1031); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1034 = $signed(_T_1032) + $signed(_T_1022); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1035 = $signed(_T_1034); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1037 = $signed(_T_1035) + $signed(_T_1023); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1038 = $signed(_T_1037); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1040 = $signed(_T_1038) + $signed(_T_1024); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1041 = $signed(_T_1040); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1043 = $signed(_T_1041) + $signed(_T_1025); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1044 = $signed(_T_1043); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1046 = $signed(_T_1044) + $signed(_T_1026); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1047 = $signed(_T_1046); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1049 = $signed(_T_1047) + $signed(_T_1027); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1050 = $signed(_T_1049); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1052 = $signed(_T_1050) + $signed(_T_1028); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1053 = $signed(_T_1052); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1055 = $signed(_T_1053) + $signed(_T_1029); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1056 = $signed(_T_1055); // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_152 = {{8{io_outputBias[31]}},io_outputBias}; // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_153 = $signed(_GEN_152) << 8; // @[FixedPointTypeClass.scala 21:58]
  assign _GEN_154 = {{24{_GEN_153[39]}},_GEN_153}; // @[FixedPointTypeClass.scala 21:58]
  assign _T_1058 = $signed(_T_1056) + $signed(_GEN_154); // @[FixedPointTypeClass.scala 21:58]
  assign linearOut = $signed(_T_1058); // @[FixedPointTypeClass.scala 21:58]
  assign _T_1059 = $signed(linearOut) > $signed(64'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign actualVotes = _T_1059 ? $signed(linearOut) : $signed(64'sh0); // @[neuralNet.scala 69:24]
  assign finalPredict = $signed(actualVotes) > $signed(64'sh0); // @[FixedPointTypeClass.scala 56:59]
  assign io_out_valid = valReg; // @[neuralNet.scala 81:16]
  assign io_out_bits = outReg; // @[neuralNet.scala 80:15]
  assign _GEN_155 = rawVotesReg[63:8]; // @[neuralNet.scala 79:15]
  assign _GEN_156 = _GEN_155[31:0]; // @[neuralNet.scala 79:15]
  assign io_rawVotes = $signed(_GEN_156); // @[neuralNet.scala 79:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  rawVotesReg = _RAND_0[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  outReg = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  valReg = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (io_in_valid) begin
      if (_T_1059) begin
        rawVotesReg <= linearOut;
      end else begin
        rawVotesReg <= 64'sh0;
      end
    end
    if (io_in_valid) begin
      outReg <= finalPredict;
    end
    valReg <= io_in_valid;
  end
endmodule
module WellnessModule(
  input         clock,
  input         reset,
  input         io_streamIn_valid,
  input  [31:0] io_streamIn_bits,
  input         io_in_valid,
  input  [31:0] io_in_bits,
  input  [31:0] io_inConf_bits_confneuralNetsinputWeights_0_0,
  input  [31:0] io_inConf_bits_confneuralNetsinputWeights_0_1,
  input  [31:0] io_inConf_bits_confneuralNetsinputWeights_0_2,
  input  [31:0] io_inConf_bits_confneuralNetsinputWeights_0_3,
  input  [31:0] io_inConf_bits_confneuralNetsinputWeights_1_0,
  input  [31:0] io_inConf_bits_confneuralNetsinputWeights_1_1,
  input  [31:0] io_inConf_bits_confneuralNetsinputWeights_1_2,
  input  [31:0] io_inConf_bits_confneuralNetsinputWeights_1_3,
  input  [31:0] io_inConf_bits_confneuralNetsinputWeights_2_0,
  input  [31:0] io_inConf_bits_confneuralNetsinputWeights_2_1,
  input  [31:0] io_inConf_bits_confneuralNetsinputWeights_2_2,
  input  [31:0] io_inConf_bits_confneuralNetsinputWeights_2_3,
  input  [31:0] io_inConf_bits_confneuralNetsinputWeights_3_0,
  input  [31:0] io_inConf_bits_confneuralNetsinputWeights_3_1,
  input  [31:0] io_inConf_bits_confneuralNetsinputWeights_3_2,
  input  [31:0] io_inConf_bits_confneuralNetsinputWeights_3_3,
  input  [31:0] io_inConf_bits_confneuralNetsinputWeights_4_0,
  input  [31:0] io_inConf_bits_confneuralNetsinputWeights_4_1,
  input  [31:0] io_inConf_bits_confneuralNetsinputWeights_4_2,
  input  [31:0] io_inConf_bits_confneuralNetsinputWeights_4_3,
  input  [31:0] io_inConf_bits_confneuralNetsinputWeights_5_0,
  input  [31:0] io_inConf_bits_confneuralNetsinputWeights_5_1,
  input  [31:0] io_inConf_bits_confneuralNetsinputWeights_5_2,
  input  [31:0] io_inConf_bits_confneuralNetsinputWeights_5_3,
  input  [31:0] io_inConf_bits_confneuralNetsinputWeights_6_0,
  input  [31:0] io_inConf_bits_confneuralNetsinputWeights_6_1,
  input  [31:0] io_inConf_bits_confneuralNetsinputWeights_6_2,
  input  [31:0] io_inConf_bits_confneuralNetsinputWeights_6_3,
  input  [31:0] io_inConf_bits_confneuralNetsinputWeights_7_0,
  input  [31:0] io_inConf_bits_confneuralNetsinputWeights_7_1,
  input  [31:0] io_inConf_bits_confneuralNetsinputWeights_7_2,
  input  [31:0] io_inConf_bits_confneuralNetsinputWeights_7_3,
  input  [31:0] io_inConf_bits_confneuralNetsinputWeights_8_0,
  input  [31:0] io_inConf_bits_confneuralNetsinputWeights_8_1,
  input  [31:0] io_inConf_bits_confneuralNetsinputWeights_8_2,
  input  [31:0] io_inConf_bits_confneuralNetsinputWeights_8_3,
  input  [31:0] io_inConf_bits_confneuralNetsinputWeights_9_0,
  input  [31:0] io_inConf_bits_confneuralNetsinputWeights_9_1,
  input  [31:0] io_inConf_bits_confneuralNetsinputWeights_9_2,
  input  [31:0] io_inConf_bits_confneuralNetsinputWeights_9_3,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_0_0,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_0_1,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_0_2,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_0_3,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_0_4,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_0_5,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_0_6,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_0_7,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_0_8,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_0_9,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_1_0,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_1_1,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_1_2,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_1_3,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_1_4,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_1_5,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_1_6,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_1_7,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_1_8,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_1_9,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_2_0,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_2_1,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_2_2,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_2_3,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_2_4,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_2_5,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_2_6,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_2_7,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_2_8,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_2_9,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_3_0,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_3_1,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_3_2,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_3_3,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_3_4,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_3_5,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_3_6,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_3_7,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_3_8,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_3_9,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_4_0,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_4_1,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_4_2,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_4_3,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_4_4,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_4_5,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_4_6,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_4_7,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_4_8,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_4_9,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_5_0,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_5_1,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_5_2,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_5_3,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_5_4,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_5_5,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_5_6,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_5_7,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_5_8,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_5_9,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_6_0,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_6_1,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_6_2,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_6_3,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_6_4,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_6_5,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_6_6,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_6_7,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_6_8,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_6_9,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_7_0,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_7_1,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_7_2,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_7_3,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_7_4,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_7_5,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_7_6,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_7_7,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_7_8,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_7_9,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_8_0,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_8_1,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_8_2,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_8_3,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_8_4,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_8_5,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_8_6,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_8_7,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_8_8,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_8_9,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_9_0,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_9_1,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_9_2,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_9_3,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_9_4,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_9_5,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_9_6,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_9_7,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_9_8,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_9_9,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_10_0,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_10_1,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_10_2,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_10_3,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_10_4,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_10_5,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_10_6,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_10_7,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_10_8,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_10_9,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_11_0,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_11_1,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_11_2,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_11_3,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_11_4,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_11_5,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_11_6,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_11_7,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_11_8,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_11_9,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_12_0,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_12_1,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_12_2,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_12_3,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_12_4,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_12_5,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_12_6,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_12_7,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_12_8,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_12_9,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_13_0,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_13_1,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_13_2,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_13_3,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_13_4,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_13_5,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_13_6,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_13_7,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_13_8,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_13_9,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_14_0,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_14_1,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_14_2,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_14_3,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_14_4,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_14_5,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_14_6,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_14_7,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_14_8,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_14_9,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_15_0,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_15_1,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_15_2,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_15_3,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_15_4,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_15_5,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_15_6,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_15_7,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_15_8,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_15_9,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_16_0,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_16_1,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_16_2,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_16_3,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_16_4,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_16_5,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_16_6,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_16_7,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_16_8,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_16_9,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_17_0,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_17_1,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_17_2,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_17_3,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_17_4,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_17_5,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_17_6,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_17_7,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_17_8,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_17_9,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_18_0,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_18_1,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_18_2,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_18_3,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_18_4,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_18_5,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_18_6,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_18_7,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_18_8,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_18_9,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_19_0,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_19_1,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_19_2,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_19_3,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_19_4,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_19_5,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_19_6,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_19_7,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_19_8,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_19_9,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_20_0,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_20_1,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_20_2,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_20_3,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_20_4,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_20_5,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_20_6,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_20_7,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_20_8,
  input  [31:0] io_inConf_bits_confneuralNetsmidAndOutputWeights_20_9,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVecs_0_0,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVecs_0_1,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVecs_0_2,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVecs_0_3,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVecs_0_4,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVecs_0_5,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVecs_0_6,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVecs_0_7,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVecs_0_8,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVecs_0_9,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVecs_1_0,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVecs_1_1,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVecs_1_2,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVecs_1_3,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVecs_1_4,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVecs_1_5,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVecs_1_6,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVecs_1_7,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVecs_1_8,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVecs_1_9,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVecs_2_0,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVecs_2_1,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVecs_2_2,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVecs_2_3,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVecs_2_4,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVecs_2_5,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVecs_2_6,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVecs_2_7,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVecs_2_8,
  input  [31:0] io_inConf_bits_confneuralNetsbiasVecs_2_9,
  input  [31:0] io_inConf_bits_confneuralNetsoutputBias_0,
  input         io_inConf_bits_confInputMuxSel,
  output        io_out_valid,
  output        io_out_bits,
  output [31:0] io_rawVotes
);
  wire  filter1_clock; // @[Wellness.scala 255:23]
  wire  filter1_reset; // @[Wellness.scala 255:23]
  wire  filter1_io_in_valid; // @[Wellness.scala 255:23]
  wire [31:0] filter1_io_in_bits; // @[Wellness.scala 255:23]
  wire  filter1_io_out_valid; // @[Wellness.scala 255:23]
  wire [31:0] filter1_io_out_bits; // @[Wellness.scala 255:23]
  wire  lineLength1_clock; // @[Wellness.scala 256:27]
  wire  lineLength1_reset; // @[Wellness.scala 256:27]
  wire  lineLength1_io_in_valid; // @[Wellness.scala 256:27]
  wire [31:0] lineLength1_io_in_bits; // @[Wellness.scala 256:27]
  wire  lineLength1_io_out_valid; // @[Wellness.scala 256:27]
  wire [31:0] lineLength1_io_out_bits; // @[Wellness.scala 256:27]
  wire  filterAlpha_clock; // @[Wellness.scala 258:27]
  wire  filterAlpha_reset; // @[Wellness.scala 258:27]
  wire  filterAlpha_io_in_valid; // @[Wellness.scala 258:27]
  wire [31:0] filterAlpha_io_in_bits; // @[Wellness.scala 258:27]
  wire  filterAlpha_io_out_valid; // @[Wellness.scala 258:27]
  wire [31:0] filterAlpha_io_out_bits; // @[Wellness.scala 258:27]
  wire  filterBeta_clock; // @[Wellness.scala 259:26]
  wire  filterBeta_reset; // @[Wellness.scala 259:26]
  wire  filterBeta_io_in_valid; // @[Wellness.scala 259:26]
  wire [31:0] filterBeta_io_in_bits; // @[Wellness.scala 259:26]
  wire  filterBeta_io_out_valid; // @[Wellness.scala 259:26]
  wire [31:0] filterBeta_io_out_bits; // @[Wellness.scala 259:26]
  wire  filterGamma_clock; // @[Wellness.scala 260:27]
  wire  filterGamma_reset; // @[Wellness.scala 260:27]
  wire  filterGamma_io_in_valid; // @[Wellness.scala 260:27]
  wire [31:0] filterGamma_io_in_bits; // @[Wellness.scala 260:27]
  wire  filterGamma_io_out_valid; // @[Wellness.scala 260:27]
  wire [31:0] filterGamma_io_out_bits; // @[Wellness.scala 260:27]
  wire  bandpowerAlpha_clock; // @[Wellness.scala 262:30]
  wire  bandpowerAlpha_reset; // @[Wellness.scala 262:30]
  wire  bandpowerAlpha_io_in_valid; // @[Wellness.scala 262:30]
  wire [31:0] bandpowerAlpha_io_in_bits; // @[Wellness.scala 262:30]
  wire  bandpowerAlpha_io_out_valid; // @[Wellness.scala 262:30]
  wire [31:0] bandpowerAlpha_io_out_bits; // @[Wellness.scala 262:30]
  wire  bandpowerBeta_clock; // @[Wellness.scala 263:29]
  wire  bandpowerBeta_reset; // @[Wellness.scala 263:29]
  wire  bandpowerBeta_io_in_valid; // @[Wellness.scala 263:29]
  wire [31:0] bandpowerBeta_io_in_bits; // @[Wellness.scala 263:29]
  wire  bandpowerBeta_io_out_valid; // @[Wellness.scala 263:29]
  wire [31:0] bandpowerBeta_io_out_bits; // @[Wellness.scala 263:29]
  wire  bandpowerGamma_clock; // @[Wellness.scala 264:30]
  wire  bandpowerGamma_reset; // @[Wellness.scala 264:30]
  wire  bandpowerGamma_io_in_valid; // @[Wellness.scala 264:30]
  wire [31:0] bandpowerGamma_io_in_bits; // @[Wellness.scala 264:30]
  wire  bandpowerGamma_io_out_valid; // @[Wellness.scala 264:30]
  wire [31:0] bandpowerGamma_io_out_bits; // @[Wellness.scala 264:30]
  wire  neuralNets_clock; // @[Wellness.scala 266:26]
  wire  neuralNets_io_in_valid; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_in_bits_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_in_bits_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_in_bits_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_in_bits_3; // @[Wellness.scala 266:26]
  wire  neuralNets_io_out_valid; // @[Wellness.scala 266:26]
  wire  neuralNets_io_out_bits; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_inputWeights_0_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_inputWeights_0_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_inputWeights_0_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_inputWeights_0_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_inputWeights_1_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_inputWeights_1_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_inputWeights_1_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_inputWeights_1_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_inputWeights_2_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_inputWeights_2_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_inputWeights_2_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_inputWeights_2_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_inputWeights_3_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_inputWeights_3_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_inputWeights_3_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_inputWeights_3_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_inputWeights_4_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_inputWeights_4_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_inputWeights_4_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_inputWeights_4_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_inputWeights_5_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_inputWeights_5_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_inputWeights_5_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_inputWeights_5_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_inputWeights_6_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_inputWeights_6_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_inputWeights_6_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_inputWeights_6_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_inputWeights_7_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_inputWeights_7_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_inputWeights_7_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_inputWeights_7_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_inputWeights_8_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_inputWeights_8_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_inputWeights_8_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_inputWeights_8_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_inputWeights_9_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_inputWeights_9_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_inputWeights_9_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_inputWeights_9_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_0_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_0_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_0_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_0_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_0_4; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_0_5; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_0_6; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_0_7; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_0_8; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_0_9; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_1_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_1_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_1_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_1_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_1_4; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_1_5; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_1_6; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_1_7; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_1_8; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_1_9; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_2_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_2_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_2_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_2_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_2_4; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_2_5; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_2_6; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_2_7; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_2_8; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_2_9; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_3_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_3_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_3_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_3_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_3_4; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_3_5; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_3_6; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_3_7; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_3_8; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_3_9; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_4_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_4_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_4_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_4_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_4_4; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_4_5; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_4_6; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_4_7; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_4_8; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_4_9; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_5_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_5_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_5_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_5_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_5_4; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_5_5; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_5_6; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_5_7; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_5_8; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_5_9; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_6_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_6_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_6_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_6_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_6_4; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_6_5; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_6_6; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_6_7; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_6_8; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_6_9; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_7_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_7_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_7_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_7_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_7_4; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_7_5; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_7_6; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_7_7; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_7_8; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_7_9; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_8_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_8_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_8_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_8_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_8_4; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_8_5; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_8_6; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_8_7; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_8_8; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_8_9; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_9_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_9_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_9_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_9_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_9_4; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_9_5; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_9_6; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_9_7; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_9_8; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_9_9; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_10_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_10_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_10_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_10_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_10_4; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_10_5; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_10_6; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_10_7; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_10_8; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_10_9; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_11_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_11_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_11_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_11_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_11_4; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_11_5; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_11_6; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_11_7; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_11_8; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_11_9; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_12_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_12_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_12_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_12_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_12_4; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_12_5; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_12_6; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_12_7; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_12_8; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_12_9; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_13_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_13_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_13_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_13_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_13_4; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_13_5; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_13_6; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_13_7; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_13_8; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_13_9; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_14_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_14_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_14_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_14_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_14_4; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_14_5; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_14_6; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_14_7; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_14_8; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_14_9; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_15_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_15_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_15_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_15_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_15_4; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_15_5; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_15_6; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_15_7; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_15_8; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_15_9; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_16_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_16_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_16_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_16_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_16_4; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_16_5; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_16_6; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_16_7; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_16_8; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_16_9; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_17_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_17_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_17_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_17_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_17_4; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_17_5; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_17_6; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_17_7; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_17_8; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_17_9; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_18_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_18_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_18_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_18_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_18_4; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_18_5; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_18_6; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_18_7; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_18_8; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_18_9; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_19_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_19_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_19_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_19_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_19_4; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_19_5; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_19_6; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_19_7; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_19_8; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_19_9; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_20_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_20_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_20_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_20_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_20_4; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_20_5; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_20_6; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_20_7; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_20_8; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_midAndOutputWeights_20_9; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVecs_0_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVecs_0_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVecs_0_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVecs_0_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVecs_0_4; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVecs_0_5; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVecs_0_6; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVecs_0_7; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVecs_0_8; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVecs_0_9; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVecs_1_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVecs_1_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVecs_1_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVecs_1_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVecs_1_4; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVecs_1_5; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVecs_1_6; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVecs_1_7; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVecs_1_8; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVecs_1_9; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVecs_2_0; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVecs_2_1; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVecs_2_2; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVecs_2_3; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVecs_2_4; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVecs_2_5; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVecs_2_6; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVecs_2_7; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVecs_2_8; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_biasVecs_2_9; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_outputBias; // @[Wellness.scala 266:26]
  wire [31:0] neuralNets_io_rawVotes; // @[Wellness.scala 266:26]
  wire [31:0] _T_1; // @[Wellness.scala 271:80]
  wire [31:0] _T_2; // @[Wellness.scala 271:80]
  wire [31:0] _T_4; // @[Wellness.scala 271:125]
  wire [31:0] _T_5; // @[Wellness.scala 271:125]
  wire [31:0] _T_10; // @[Wellness.scala 283:57]
  wire [31:0] _T_22; // @[Wellness.scala 314:65]
  reg [31:0] lineLength1Reg1; // @[Wellness.scala 314:32]
  reg [31:0] _RAND_0;
  reg  lineLength1Valid1; // @[Wellness.scala 316:34]
  reg [31:0] _RAND_1;
  wire [31:0] _T_25; // @[Wellness.scala 327:58]
  wire [31:0] _T_28; // @[Wellness.scala 328:57]
  wire [31:0] _T_31; // @[Wellness.scala 329:58]
  wire [31:0] _T_34; // @[Wellness.scala 330:47]
  wire  _T_36; // @[Wellness.scala 332:48]
  wire  _T_37; // @[Wellness.scala 332:79]
  ConstantCoefficientFIRFilter filter1 ( // @[Wellness.scala 255:23]
    .clock(filter1_clock),
    .reset(filter1_reset),
    .io_in_valid(filter1_io_in_valid),
    .io_in_bits(filter1_io_in_bits),
    .io_out_valid(filter1_io_out_valid),
    .io_out_bits(filter1_io_out_bits)
  );
  lineLength lineLength1 ( // @[Wellness.scala 256:27]
    .clock(lineLength1_clock),
    .reset(lineLength1_reset),
    .io_in_valid(lineLength1_io_in_valid),
    .io_in_bits(lineLength1_io_in_bits),
    .io_out_valid(lineLength1_io_out_valid),
    .io_out_bits(lineLength1_io_out_bits)
  );
  ConstantCoefficientFIRFilter filterAlpha ( // @[Wellness.scala 258:27]
    .clock(filterAlpha_clock),
    .reset(filterAlpha_reset),
    .io_in_valid(filterAlpha_io_in_valid),
    .io_in_bits(filterAlpha_io_in_bits),
    .io_out_valid(filterAlpha_io_out_valid),
    .io_out_bits(filterAlpha_io_out_bits)
  );
  ConstantCoefficientFIRFilter filterBeta ( // @[Wellness.scala 259:26]
    .clock(filterBeta_clock),
    .reset(filterBeta_reset),
    .io_in_valid(filterBeta_io_in_valid),
    .io_in_bits(filterBeta_io_in_bits),
    .io_out_valid(filterBeta_io_out_valid),
    .io_out_bits(filterBeta_io_out_bits)
  );
  ConstantCoefficientFIRFilter filterGamma ( // @[Wellness.scala 260:27]
    .clock(filterGamma_clock),
    .reset(filterGamma_reset),
    .io_in_valid(filterGamma_io_in_valid),
    .io_in_bits(filterGamma_io_in_bits),
    .io_out_valid(filterGamma_io_out_valid),
    .io_out_bits(filterGamma_io_out_bits)
  );
  sumSquares bandpowerAlpha ( // @[Wellness.scala 262:30]
    .clock(bandpowerAlpha_clock),
    .reset(bandpowerAlpha_reset),
    .io_in_valid(bandpowerAlpha_io_in_valid),
    .io_in_bits(bandpowerAlpha_io_in_bits),
    .io_out_valid(bandpowerAlpha_io_out_valid),
    .io_out_bits(bandpowerAlpha_io_out_bits)
  );
  sumSquares bandpowerBeta ( // @[Wellness.scala 263:29]
    .clock(bandpowerBeta_clock),
    .reset(bandpowerBeta_reset),
    .io_in_valid(bandpowerBeta_io_in_valid),
    .io_in_bits(bandpowerBeta_io_in_bits),
    .io_out_valid(bandpowerBeta_io_out_valid),
    .io_out_bits(bandpowerBeta_io_out_bits)
  );
  sumSquares bandpowerGamma ( // @[Wellness.scala 264:30]
    .clock(bandpowerGamma_clock),
    .reset(bandpowerGamma_reset),
    .io_in_valid(bandpowerGamma_io_in_valid),
    .io_in_bits(bandpowerGamma_io_in_bits),
    .io_out_valid(bandpowerGamma_io_out_valid),
    .io_out_bits(bandpowerGamma_io_out_bits)
  );
  NeuralNet neuralNets ( // @[Wellness.scala 266:26]
    .clock(neuralNets_clock),
    .io_in_valid(neuralNets_io_in_valid),
    .io_in_bits_0(neuralNets_io_in_bits_0),
    .io_in_bits_1(neuralNets_io_in_bits_1),
    .io_in_bits_2(neuralNets_io_in_bits_2),
    .io_in_bits_3(neuralNets_io_in_bits_3),
    .io_out_valid(neuralNets_io_out_valid),
    .io_out_bits(neuralNets_io_out_bits),
    .io_inputWeights_0_0(neuralNets_io_inputWeights_0_0),
    .io_inputWeights_0_1(neuralNets_io_inputWeights_0_1),
    .io_inputWeights_0_2(neuralNets_io_inputWeights_0_2),
    .io_inputWeights_0_3(neuralNets_io_inputWeights_0_3),
    .io_inputWeights_1_0(neuralNets_io_inputWeights_1_0),
    .io_inputWeights_1_1(neuralNets_io_inputWeights_1_1),
    .io_inputWeights_1_2(neuralNets_io_inputWeights_1_2),
    .io_inputWeights_1_3(neuralNets_io_inputWeights_1_3),
    .io_inputWeights_2_0(neuralNets_io_inputWeights_2_0),
    .io_inputWeights_2_1(neuralNets_io_inputWeights_2_1),
    .io_inputWeights_2_2(neuralNets_io_inputWeights_2_2),
    .io_inputWeights_2_3(neuralNets_io_inputWeights_2_3),
    .io_inputWeights_3_0(neuralNets_io_inputWeights_3_0),
    .io_inputWeights_3_1(neuralNets_io_inputWeights_3_1),
    .io_inputWeights_3_2(neuralNets_io_inputWeights_3_2),
    .io_inputWeights_3_3(neuralNets_io_inputWeights_3_3),
    .io_inputWeights_4_0(neuralNets_io_inputWeights_4_0),
    .io_inputWeights_4_1(neuralNets_io_inputWeights_4_1),
    .io_inputWeights_4_2(neuralNets_io_inputWeights_4_2),
    .io_inputWeights_4_3(neuralNets_io_inputWeights_4_3),
    .io_inputWeights_5_0(neuralNets_io_inputWeights_5_0),
    .io_inputWeights_5_1(neuralNets_io_inputWeights_5_1),
    .io_inputWeights_5_2(neuralNets_io_inputWeights_5_2),
    .io_inputWeights_5_3(neuralNets_io_inputWeights_5_3),
    .io_inputWeights_6_0(neuralNets_io_inputWeights_6_0),
    .io_inputWeights_6_1(neuralNets_io_inputWeights_6_1),
    .io_inputWeights_6_2(neuralNets_io_inputWeights_6_2),
    .io_inputWeights_6_3(neuralNets_io_inputWeights_6_3),
    .io_inputWeights_7_0(neuralNets_io_inputWeights_7_0),
    .io_inputWeights_7_1(neuralNets_io_inputWeights_7_1),
    .io_inputWeights_7_2(neuralNets_io_inputWeights_7_2),
    .io_inputWeights_7_3(neuralNets_io_inputWeights_7_3),
    .io_inputWeights_8_0(neuralNets_io_inputWeights_8_0),
    .io_inputWeights_8_1(neuralNets_io_inputWeights_8_1),
    .io_inputWeights_8_2(neuralNets_io_inputWeights_8_2),
    .io_inputWeights_8_3(neuralNets_io_inputWeights_8_3),
    .io_inputWeights_9_0(neuralNets_io_inputWeights_9_0),
    .io_inputWeights_9_1(neuralNets_io_inputWeights_9_1),
    .io_inputWeights_9_2(neuralNets_io_inputWeights_9_2),
    .io_inputWeights_9_3(neuralNets_io_inputWeights_9_3),
    .io_midAndOutputWeights_0_0(neuralNets_io_midAndOutputWeights_0_0),
    .io_midAndOutputWeights_0_1(neuralNets_io_midAndOutputWeights_0_1),
    .io_midAndOutputWeights_0_2(neuralNets_io_midAndOutputWeights_0_2),
    .io_midAndOutputWeights_0_3(neuralNets_io_midAndOutputWeights_0_3),
    .io_midAndOutputWeights_0_4(neuralNets_io_midAndOutputWeights_0_4),
    .io_midAndOutputWeights_0_5(neuralNets_io_midAndOutputWeights_0_5),
    .io_midAndOutputWeights_0_6(neuralNets_io_midAndOutputWeights_0_6),
    .io_midAndOutputWeights_0_7(neuralNets_io_midAndOutputWeights_0_7),
    .io_midAndOutputWeights_0_8(neuralNets_io_midAndOutputWeights_0_8),
    .io_midAndOutputWeights_0_9(neuralNets_io_midAndOutputWeights_0_9),
    .io_midAndOutputWeights_1_0(neuralNets_io_midAndOutputWeights_1_0),
    .io_midAndOutputWeights_1_1(neuralNets_io_midAndOutputWeights_1_1),
    .io_midAndOutputWeights_1_2(neuralNets_io_midAndOutputWeights_1_2),
    .io_midAndOutputWeights_1_3(neuralNets_io_midAndOutputWeights_1_3),
    .io_midAndOutputWeights_1_4(neuralNets_io_midAndOutputWeights_1_4),
    .io_midAndOutputWeights_1_5(neuralNets_io_midAndOutputWeights_1_5),
    .io_midAndOutputWeights_1_6(neuralNets_io_midAndOutputWeights_1_6),
    .io_midAndOutputWeights_1_7(neuralNets_io_midAndOutputWeights_1_7),
    .io_midAndOutputWeights_1_8(neuralNets_io_midAndOutputWeights_1_8),
    .io_midAndOutputWeights_1_9(neuralNets_io_midAndOutputWeights_1_9),
    .io_midAndOutputWeights_2_0(neuralNets_io_midAndOutputWeights_2_0),
    .io_midAndOutputWeights_2_1(neuralNets_io_midAndOutputWeights_2_1),
    .io_midAndOutputWeights_2_2(neuralNets_io_midAndOutputWeights_2_2),
    .io_midAndOutputWeights_2_3(neuralNets_io_midAndOutputWeights_2_3),
    .io_midAndOutputWeights_2_4(neuralNets_io_midAndOutputWeights_2_4),
    .io_midAndOutputWeights_2_5(neuralNets_io_midAndOutputWeights_2_5),
    .io_midAndOutputWeights_2_6(neuralNets_io_midAndOutputWeights_2_6),
    .io_midAndOutputWeights_2_7(neuralNets_io_midAndOutputWeights_2_7),
    .io_midAndOutputWeights_2_8(neuralNets_io_midAndOutputWeights_2_8),
    .io_midAndOutputWeights_2_9(neuralNets_io_midAndOutputWeights_2_9),
    .io_midAndOutputWeights_3_0(neuralNets_io_midAndOutputWeights_3_0),
    .io_midAndOutputWeights_3_1(neuralNets_io_midAndOutputWeights_3_1),
    .io_midAndOutputWeights_3_2(neuralNets_io_midAndOutputWeights_3_2),
    .io_midAndOutputWeights_3_3(neuralNets_io_midAndOutputWeights_3_3),
    .io_midAndOutputWeights_3_4(neuralNets_io_midAndOutputWeights_3_4),
    .io_midAndOutputWeights_3_5(neuralNets_io_midAndOutputWeights_3_5),
    .io_midAndOutputWeights_3_6(neuralNets_io_midAndOutputWeights_3_6),
    .io_midAndOutputWeights_3_7(neuralNets_io_midAndOutputWeights_3_7),
    .io_midAndOutputWeights_3_8(neuralNets_io_midAndOutputWeights_3_8),
    .io_midAndOutputWeights_3_9(neuralNets_io_midAndOutputWeights_3_9),
    .io_midAndOutputWeights_4_0(neuralNets_io_midAndOutputWeights_4_0),
    .io_midAndOutputWeights_4_1(neuralNets_io_midAndOutputWeights_4_1),
    .io_midAndOutputWeights_4_2(neuralNets_io_midAndOutputWeights_4_2),
    .io_midAndOutputWeights_4_3(neuralNets_io_midAndOutputWeights_4_3),
    .io_midAndOutputWeights_4_4(neuralNets_io_midAndOutputWeights_4_4),
    .io_midAndOutputWeights_4_5(neuralNets_io_midAndOutputWeights_4_5),
    .io_midAndOutputWeights_4_6(neuralNets_io_midAndOutputWeights_4_6),
    .io_midAndOutputWeights_4_7(neuralNets_io_midAndOutputWeights_4_7),
    .io_midAndOutputWeights_4_8(neuralNets_io_midAndOutputWeights_4_8),
    .io_midAndOutputWeights_4_9(neuralNets_io_midAndOutputWeights_4_9),
    .io_midAndOutputWeights_5_0(neuralNets_io_midAndOutputWeights_5_0),
    .io_midAndOutputWeights_5_1(neuralNets_io_midAndOutputWeights_5_1),
    .io_midAndOutputWeights_5_2(neuralNets_io_midAndOutputWeights_5_2),
    .io_midAndOutputWeights_5_3(neuralNets_io_midAndOutputWeights_5_3),
    .io_midAndOutputWeights_5_4(neuralNets_io_midAndOutputWeights_5_4),
    .io_midAndOutputWeights_5_5(neuralNets_io_midAndOutputWeights_5_5),
    .io_midAndOutputWeights_5_6(neuralNets_io_midAndOutputWeights_5_6),
    .io_midAndOutputWeights_5_7(neuralNets_io_midAndOutputWeights_5_7),
    .io_midAndOutputWeights_5_8(neuralNets_io_midAndOutputWeights_5_8),
    .io_midAndOutputWeights_5_9(neuralNets_io_midAndOutputWeights_5_9),
    .io_midAndOutputWeights_6_0(neuralNets_io_midAndOutputWeights_6_0),
    .io_midAndOutputWeights_6_1(neuralNets_io_midAndOutputWeights_6_1),
    .io_midAndOutputWeights_6_2(neuralNets_io_midAndOutputWeights_6_2),
    .io_midAndOutputWeights_6_3(neuralNets_io_midAndOutputWeights_6_3),
    .io_midAndOutputWeights_6_4(neuralNets_io_midAndOutputWeights_6_4),
    .io_midAndOutputWeights_6_5(neuralNets_io_midAndOutputWeights_6_5),
    .io_midAndOutputWeights_6_6(neuralNets_io_midAndOutputWeights_6_6),
    .io_midAndOutputWeights_6_7(neuralNets_io_midAndOutputWeights_6_7),
    .io_midAndOutputWeights_6_8(neuralNets_io_midAndOutputWeights_6_8),
    .io_midAndOutputWeights_6_9(neuralNets_io_midAndOutputWeights_6_9),
    .io_midAndOutputWeights_7_0(neuralNets_io_midAndOutputWeights_7_0),
    .io_midAndOutputWeights_7_1(neuralNets_io_midAndOutputWeights_7_1),
    .io_midAndOutputWeights_7_2(neuralNets_io_midAndOutputWeights_7_2),
    .io_midAndOutputWeights_7_3(neuralNets_io_midAndOutputWeights_7_3),
    .io_midAndOutputWeights_7_4(neuralNets_io_midAndOutputWeights_7_4),
    .io_midAndOutputWeights_7_5(neuralNets_io_midAndOutputWeights_7_5),
    .io_midAndOutputWeights_7_6(neuralNets_io_midAndOutputWeights_7_6),
    .io_midAndOutputWeights_7_7(neuralNets_io_midAndOutputWeights_7_7),
    .io_midAndOutputWeights_7_8(neuralNets_io_midAndOutputWeights_7_8),
    .io_midAndOutputWeights_7_9(neuralNets_io_midAndOutputWeights_7_9),
    .io_midAndOutputWeights_8_0(neuralNets_io_midAndOutputWeights_8_0),
    .io_midAndOutputWeights_8_1(neuralNets_io_midAndOutputWeights_8_1),
    .io_midAndOutputWeights_8_2(neuralNets_io_midAndOutputWeights_8_2),
    .io_midAndOutputWeights_8_3(neuralNets_io_midAndOutputWeights_8_3),
    .io_midAndOutputWeights_8_4(neuralNets_io_midAndOutputWeights_8_4),
    .io_midAndOutputWeights_8_5(neuralNets_io_midAndOutputWeights_8_5),
    .io_midAndOutputWeights_8_6(neuralNets_io_midAndOutputWeights_8_6),
    .io_midAndOutputWeights_8_7(neuralNets_io_midAndOutputWeights_8_7),
    .io_midAndOutputWeights_8_8(neuralNets_io_midAndOutputWeights_8_8),
    .io_midAndOutputWeights_8_9(neuralNets_io_midAndOutputWeights_8_9),
    .io_midAndOutputWeights_9_0(neuralNets_io_midAndOutputWeights_9_0),
    .io_midAndOutputWeights_9_1(neuralNets_io_midAndOutputWeights_9_1),
    .io_midAndOutputWeights_9_2(neuralNets_io_midAndOutputWeights_9_2),
    .io_midAndOutputWeights_9_3(neuralNets_io_midAndOutputWeights_9_3),
    .io_midAndOutputWeights_9_4(neuralNets_io_midAndOutputWeights_9_4),
    .io_midAndOutputWeights_9_5(neuralNets_io_midAndOutputWeights_9_5),
    .io_midAndOutputWeights_9_6(neuralNets_io_midAndOutputWeights_9_6),
    .io_midAndOutputWeights_9_7(neuralNets_io_midAndOutputWeights_9_7),
    .io_midAndOutputWeights_9_8(neuralNets_io_midAndOutputWeights_9_8),
    .io_midAndOutputWeights_9_9(neuralNets_io_midAndOutputWeights_9_9),
    .io_midAndOutputWeights_10_0(neuralNets_io_midAndOutputWeights_10_0),
    .io_midAndOutputWeights_10_1(neuralNets_io_midAndOutputWeights_10_1),
    .io_midAndOutputWeights_10_2(neuralNets_io_midAndOutputWeights_10_2),
    .io_midAndOutputWeights_10_3(neuralNets_io_midAndOutputWeights_10_3),
    .io_midAndOutputWeights_10_4(neuralNets_io_midAndOutputWeights_10_4),
    .io_midAndOutputWeights_10_5(neuralNets_io_midAndOutputWeights_10_5),
    .io_midAndOutputWeights_10_6(neuralNets_io_midAndOutputWeights_10_6),
    .io_midAndOutputWeights_10_7(neuralNets_io_midAndOutputWeights_10_7),
    .io_midAndOutputWeights_10_8(neuralNets_io_midAndOutputWeights_10_8),
    .io_midAndOutputWeights_10_9(neuralNets_io_midAndOutputWeights_10_9),
    .io_midAndOutputWeights_11_0(neuralNets_io_midAndOutputWeights_11_0),
    .io_midAndOutputWeights_11_1(neuralNets_io_midAndOutputWeights_11_1),
    .io_midAndOutputWeights_11_2(neuralNets_io_midAndOutputWeights_11_2),
    .io_midAndOutputWeights_11_3(neuralNets_io_midAndOutputWeights_11_3),
    .io_midAndOutputWeights_11_4(neuralNets_io_midAndOutputWeights_11_4),
    .io_midAndOutputWeights_11_5(neuralNets_io_midAndOutputWeights_11_5),
    .io_midAndOutputWeights_11_6(neuralNets_io_midAndOutputWeights_11_6),
    .io_midAndOutputWeights_11_7(neuralNets_io_midAndOutputWeights_11_7),
    .io_midAndOutputWeights_11_8(neuralNets_io_midAndOutputWeights_11_8),
    .io_midAndOutputWeights_11_9(neuralNets_io_midAndOutputWeights_11_9),
    .io_midAndOutputWeights_12_0(neuralNets_io_midAndOutputWeights_12_0),
    .io_midAndOutputWeights_12_1(neuralNets_io_midAndOutputWeights_12_1),
    .io_midAndOutputWeights_12_2(neuralNets_io_midAndOutputWeights_12_2),
    .io_midAndOutputWeights_12_3(neuralNets_io_midAndOutputWeights_12_3),
    .io_midAndOutputWeights_12_4(neuralNets_io_midAndOutputWeights_12_4),
    .io_midAndOutputWeights_12_5(neuralNets_io_midAndOutputWeights_12_5),
    .io_midAndOutputWeights_12_6(neuralNets_io_midAndOutputWeights_12_6),
    .io_midAndOutputWeights_12_7(neuralNets_io_midAndOutputWeights_12_7),
    .io_midAndOutputWeights_12_8(neuralNets_io_midAndOutputWeights_12_8),
    .io_midAndOutputWeights_12_9(neuralNets_io_midAndOutputWeights_12_9),
    .io_midAndOutputWeights_13_0(neuralNets_io_midAndOutputWeights_13_0),
    .io_midAndOutputWeights_13_1(neuralNets_io_midAndOutputWeights_13_1),
    .io_midAndOutputWeights_13_2(neuralNets_io_midAndOutputWeights_13_2),
    .io_midAndOutputWeights_13_3(neuralNets_io_midAndOutputWeights_13_3),
    .io_midAndOutputWeights_13_4(neuralNets_io_midAndOutputWeights_13_4),
    .io_midAndOutputWeights_13_5(neuralNets_io_midAndOutputWeights_13_5),
    .io_midAndOutputWeights_13_6(neuralNets_io_midAndOutputWeights_13_6),
    .io_midAndOutputWeights_13_7(neuralNets_io_midAndOutputWeights_13_7),
    .io_midAndOutputWeights_13_8(neuralNets_io_midAndOutputWeights_13_8),
    .io_midAndOutputWeights_13_9(neuralNets_io_midAndOutputWeights_13_9),
    .io_midAndOutputWeights_14_0(neuralNets_io_midAndOutputWeights_14_0),
    .io_midAndOutputWeights_14_1(neuralNets_io_midAndOutputWeights_14_1),
    .io_midAndOutputWeights_14_2(neuralNets_io_midAndOutputWeights_14_2),
    .io_midAndOutputWeights_14_3(neuralNets_io_midAndOutputWeights_14_3),
    .io_midAndOutputWeights_14_4(neuralNets_io_midAndOutputWeights_14_4),
    .io_midAndOutputWeights_14_5(neuralNets_io_midAndOutputWeights_14_5),
    .io_midAndOutputWeights_14_6(neuralNets_io_midAndOutputWeights_14_6),
    .io_midAndOutputWeights_14_7(neuralNets_io_midAndOutputWeights_14_7),
    .io_midAndOutputWeights_14_8(neuralNets_io_midAndOutputWeights_14_8),
    .io_midAndOutputWeights_14_9(neuralNets_io_midAndOutputWeights_14_9),
    .io_midAndOutputWeights_15_0(neuralNets_io_midAndOutputWeights_15_0),
    .io_midAndOutputWeights_15_1(neuralNets_io_midAndOutputWeights_15_1),
    .io_midAndOutputWeights_15_2(neuralNets_io_midAndOutputWeights_15_2),
    .io_midAndOutputWeights_15_3(neuralNets_io_midAndOutputWeights_15_3),
    .io_midAndOutputWeights_15_4(neuralNets_io_midAndOutputWeights_15_4),
    .io_midAndOutputWeights_15_5(neuralNets_io_midAndOutputWeights_15_5),
    .io_midAndOutputWeights_15_6(neuralNets_io_midAndOutputWeights_15_6),
    .io_midAndOutputWeights_15_7(neuralNets_io_midAndOutputWeights_15_7),
    .io_midAndOutputWeights_15_8(neuralNets_io_midAndOutputWeights_15_8),
    .io_midAndOutputWeights_15_9(neuralNets_io_midAndOutputWeights_15_9),
    .io_midAndOutputWeights_16_0(neuralNets_io_midAndOutputWeights_16_0),
    .io_midAndOutputWeights_16_1(neuralNets_io_midAndOutputWeights_16_1),
    .io_midAndOutputWeights_16_2(neuralNets_io_midAndOutputWeights_16_2),
    .io_midAndOutputWeights_16_3(neuralNets_io_midAndOutputWeights_16_3),
    .io_midAndOutputWeights_16_4(neuralNets_io_midAndOutputWeights_16_4),
    .io_midAndOutputWeights_16_5(neuralNets_io_midAndOutputWeights_16_5),
    .io_midAndOutputWeights_16_6(neuralNets_io_midAndOutputWeights_16_6),
    .io_midAndOutputWeights_16_7(neuralNets_io_midAndOutputWeights_16_7),
    .io_midAndOutputWeights_16_8(neuralNets_io_midAndOutputWeights_16_8),
    .io_midAndOutputWeights_16_9(neuralNets_io_midAndOutputWeights_16_9),
    .io_midAndOutputWeights_17_0(neuralNets_io_midAndOutputWeights_17_0),
    .io_midAndOutputWeights_17_1(neuralNets_io_midAndOutputWeights_17_1),
    .io_midAndOutputWeights_17_2(neuralNets_io_midAndOutputWeights_17_2),
    .io_midAndOutputWeights_17_3(neuralNets_io_midAndOutputWeights_17_3),
    .io_midAndOutputWeights_17_4(neuralNets_io_midAndOutputWeights_17_4),
    .io_midAndOutputWeights_17_5(neuralNets_io_midAndOutputWeights_17_5),
    .io_midAndOutputWeights_17_6(neuralNets_io_midAndOutputWeights_17_6),
    .io_midAndOutputWeights_17_7(neuralNets_io_midAndOutputWeights_17_7),
    .io_midAndOutputWeights_17_8(neuralNets_io_midAndOutputWeights_17_8),
    .io_midAndOutputWeights_17_9(neuralNets_io_midAndOutputWeights_17_9),
    .io_midAndOutputWeights_18_0(neuralNets_io_midAndOutputWeights_18_0),
    .io_midAndOutputWeights_18_1(neuralNets_io_midAndOutputWeights_18_1),
    .io_midAndOutputWeights_18_2(neuralNets_io_midAndOutputWeights_18_2),
    .io_midAndOutputWeights_18_3(neuralNets_io_midAndOutputWeights_18_3),
    .io_midAndOutputWeights_18_4(neuralNets_io_midAndOutputWeights_18_4),
    .io_midAndOutputWeights_18_5(neuralNets_io_midAndOutputWeights_18_5),
    .io_midAndOutputWeights_18_6(neuralNets_io_midAndOutputWeights_18_6),
    .io_midAndOutputWeights_18_7(neuralNets_io_midAndOutputWeights_18_7),
    .io_midAndOutputWeights_18_8(neuralNets_io_midAndOutputWeights_18_8),
    .io_midAndOutputWeights_18_9(neuralNets_io_midAndOutputWeights_18_9),
    .io_midAndOutputWeights_19_0(neuralNets_io_midAndOutputWeights_19_0),
    .io_midAndOutputWeights_19_1(neuralNets_io_midAndOutputWeights_19_1),
    .io_midAndOutputWeights_19_2(neuralNets_io_midAndOutputWeights_19_2),
    .io_midAndOutputWeights_19_3(neuralNets_io_midAndOutputWeights_19_3),
    .io_midAndOutputWeights_19_4(neuralNets_io_midAndOutputWeights_19_4),
    .io_midAndOutputWeights_19_5(neuralNets_io_midAndOutputWeights_19_5),
    .io_midAndOutputWeights_19_6(neuralNets_io_midAndOutputWeights_19_6),
    .io_midAndOutputWeights_19_7(neuralNets_io_midAndOutputWeights_19_7),
    .io_midAndOutputWeights_19_8(neuralNets_io_midAndOutputWeights_19_8),
    .io_midAndOutputWeights_19_9(neuralNets_io_midAndOutputWeights_19_9),
    .io_midAndOutputWeights_20_0(neuralNets_io_midAndOutputWeights_20_0),
    .io_midAndOutputWeights_20_1(neuralNets_io_midAndOutputWeights_20_1),
    .io_midAndOutputWeights_20_2(neuralNets_io_midAndOutputWeights_20_2),
    .io_midAndOutputWeights_20_3(neuralNets_io_midAndOutputWeights_20_3),
    .io_midAndOutputWeights_20_4(neuralNets_io_midAndOutputWeights_20_4),
    .io_midAndOutputWeights_20_5(neuralNets_io_midAndOutputWeights_20_5),
    .io_midAndOutputWeights_20_6(neuralNets_io_midAndOutputWeights_20_6),
    .io_midAndOutputWeights_20_7(neuralNets_io_midAndOutputWeights_20_7),
    .io_midAndOutputWeights_20_8(neuralNets_io_midAndOutputWeights_20_8),
    .io_midAndOutputWeights_20_9(neuralNets_io_midAndOutputWeights_20_9),
    .io_biasVecs_0_0(neuralNets_io_biasVecs_0_0),
    .io_biasVecs_0_1(neuralNets_io_biasVecs_0_1),
    .io_biasVecs_0_2(neuralNets_io_biasVecs_0_2),
    .io_biasVecs_0_3(neuralNets_io_biasVecs_0_3),
    .io_biasVecs_0_4(neuralNets_io_biasVecs_0_4),
    .io_biasVecs_0_5(neuralNets_io_biasVecs_0_5),
    .io_biasVecs_0_6(neuralNets_io_biasVecs_0_6),
    .io_biasVecs_0_7(neuralNets_io_biasVecs_0_7),
    .io_biasVecs_0_8(neuralNets_io_biasVecs_0_8),
    .io_biasVecs_0_9(neuralNets_io_biasVecs_0_9),
    .io_biasVecs_1_0(neuralNets_io_biasVecs_1_0),
    .io_biasVecs_1_1(neuralNets_io_biasVecs_1_1),
    .io_biasVecs_1_2(neuralNets_io_biasVecs_1_2),
    .io_biasVecs_1_3(neuralNets_io_biasVecs_1_3),
    .io_biasVecs_1_4(neuralNets_io_biasVecs_1_4),
    .io_biasVecs_1_5(neuralNets_io_biasVecs_1_5),
    .io_biasVecs_1_6(neuralNets_io_biasVecs_1_6),
    .io_biasVecs_1_7(neuralNets_io_biasVecs_1_7),
    .io_biasVecs_1_8(neuralNets_io_biasVecs_1_8),
    .io_biasVecs_1_9(neuralNets_io_biasVecs_1_9),
    .io_biasVecs_2_0(neuralNets_io_biasVecs_2_0),
    .io_biasVecs_2_1(neuralNets_io_biasVecs_2_1),
    .io_biasVecs_2_2(neuralNets_io_biasVecs_2_2),
    .io_biasVecs_2_3(neuralNets_io_biasVecs_2_3),
    .io_biasVecs_2_4(neuralNets_io_biasVecs_2_4),
    .io_biasVecs_2_5(neuralNets_io_biasVecs_2_5),
    .io_biasVecs_2_6(neuralNets_io_biasVecs_2_6),
    .io_biasVecs_2_7(neuralNets_io_biasVecs_2_7),
    .io_biasVecs_2_8(neuralNets_io_biasVecs_2_8),
    .io_biasVecs_2_9(neuralNets_io_biasVecs_2_9),
    .io_outputBias(neuralNets_io_outputBias),
    .io_rawVotes(neuralNets_io_rawVotes)
  );
  assign _T_1 = $unsigned(io_streamIn_bits); // @[Wellness.scala 271:80]
  assign _T_2 = $signed(_T_1); // @[Wellness.scala 271:80]
  assign _T_4 = $unsigned(io_in_bits); // @[Wellness.scala 271:125]
  assign _T_5 = $signed(_T_4); // @[Wellness.scala 271:125]
  assign _T_10 = $unsigned(filter1_io_out_bits); // @[Wellness.scala 283:57]
  assign _T_22 = $unsigned(lineLength1_io_out_bits); // @[Wellness.scala 314:65]
  assign _T_25 = $unsigned(bandpowerAlpha_io_out_bits); // @[Wellness.scala 327:58]
  assign _T_28 = $unsigned(bandpowerBeta_io_out_bits); // @[Wellness.scala 328:57]
  assign _T_31 = $unsigned(bandpowerGamma_io_out_bits); // @[Wellness.scala 329:58]
  assign _T_34 = $unsigned(lineLength1Reg1); // @[Wellness.scala 330:47]
  assign _T_36 = lineLength1Valid1 & bandpowerAlpha_io_out_valid; // @[Wellness.scala 332:48]
  assign _T_37 = _T_36 & bandpowerBeta_io_out_valid; // @[Wellness.scala 332:79]
  assign io_out_valid = neuralNets_io_out_valid; // @[Wellness.scala 342:16]
  assign io_out_bits = neuralNets_io_out_bits; // @[Wellness.scala 344:15]
  assign io_rawVotes = neuralNets_io_rawVotes; // @[Wellness.scala 345:15]
  assign filter1_clock = clock;
  assign filter1_reset = reset;
  assign filter1_io_in_valid = io_inConf_bits_confInputMuxSel ? io_streamIn_valid : io_in_valid; // @[Wellness.scala 276:23]
  assign filter1_io_in_bits = io_inConf_bits_confInputMuxSel ? $signed(_T_2) : $signed(_T_5); // @[Wellness.scala 278:22]
  assign lineLength1_clock = clock;
  assign lineLength1_reset = reset;
  assign lineLength1_io_in_valid = filter1_io_out_valid; // @[Wellness.scala 281:27]
  assign lineLength1_io_in_bits = $signed(_T_10); // @[Wellness.scala 283:26]
  assign filterAlpha_clock = clock;
  assign filterAlpha_reset = reset;
  assign filterAlpha_io_in_valid = filter1_io_out_valid; // @[Wellness.scala 286:27]
  assign filterAlpha_io_in_bits = $signed(_T_10); // @[Wellness.scala 288:26]
  assign filterBeta_clock = clock;
  assign filterBeta_reset = reset;
  assign filterBeta_io_in_valid = filter1_io_out_valid; // @[Wellness.scala 290:26]
  assign filterBeta_io_in_bits = $signed(_T_10); // @[Wellness.scala 292:25]
  assign filterGamma_clock = clock;
  assign filterGamma_reset = reset;
  assign filterGamma_io_in_valid = filter1_io_out_valid; // @[Wellness.scala 294:27]
  assign filterGamma_io_in_bits = $signed(_T_10); // @[Wellness.scala 296:26]
  assign bandpowerAlpha_clock = clock;
  assign bandpowerAlpha_reset = reset;
  assign bandpowerAlpha_io_in_valid = filterAlpha_io_out_valid; // @[Wellness.scala 300:30]
  assign bandpowerAlpha_io_in_bits = filterAlpha_io_out_bits; // @[Wellness.scala 302:29]
  assign bandpowerBeta_clock = clock;
  assign bandpowerBeta_reset = reset;
  assign bandpowerBeta_io_in_valid = filterBeta_io_out_valid; // @[Wellness.scala 304:29]
  assign bandpowerBeta_io_in_bits = filterBeta_io_out_bits; // @[Wellness.scala 306:28]
  assign bandpowerGamma_clock = clock;
  assign bandpowerGamma_reset = reset;
  assign bandpowerGamma_io_in_valid = filterGamma_io_out_valid; // @[Wellness.scala 308:30]
  assign bandpowerGamma_io_in_bits = filterGamma_io_out_bits; // @[Wellness.scala 310:29]
  assign neuralNets_clock = clock;
  assign neuralNets_io_in_valid = _T_37 & bandpowerGamma_io_out_valid; // @[Wellness.scala 332:26]
  assign neuralNets_io_in_bits_0 = $signed(_T_25); // @[Wellness.scala 333:25]
  assign neuralNets_io_in_bits_1 = $signed(_T_28); // @[Wellness.scala 333:25]
  assign neuralNets_io_in_bits_2 = $signed(_T_31); // @[Wellness.scala 333:25]
  assign neuralNets_io_in_bits_3 = $signed(_T_34); // @[Wellness.scala 333:25]
  assign neuralNets_io_inputWeights_0_0 = io_inConf_bits_confneuralNetsinputWeights_0_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_inputWeights_0_1 = io_inConf_bits_confneuralNetsinputWeights_0_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_inputWeights_0_2 = io_inConf_bits_confneuralNetsinputWeights_0_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_inputWeights_0_3 = io_inConf_bits_confneuralNetsinputWeights_0_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_inputWeights_1_0 = io_inConf_bits_confneuralNetsinputWeights_1_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_inputWeights_1_1 = io_inConf_bits_confneuralNetsinputWeights_1_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_inputWeights_1_2 = io_inConf_bits_confneuralNetsinputWeights_1_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_inputWeights_1_3 = io_inConf_bits_confneuralNetsinputWeights_1_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_inputWeights_2_0 = io_inConf_bits_confneuralNetsinputWeights_2_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_inputWeights_2_1 = io_inConf_bits_confneuralNetsinputWeights_2_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_inputWeights_2_2 = io_inConf_bits_confneuralNetsinputWeights_2_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_inputWeights_2_3 = io_inConf_bits_confneuralNetsinputWeights_2_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_inputWeights_3_0 = io_inConf_bits_confneuralNetsinputWeights_3_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_inputWeights_3_1 = io_inConf_bits_confneuralNetsinputWeights_3_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_inputWeights_3_2 = io_inConf_bits_confneuralNetsinputWeights_3_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_inputWeights_3_3 = io_inConf_bits_confneuralNetsinputWeights_3_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_inputWeights_4_0 = io_inConf_bits_confneuralNetsinputWeights_4_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_inputWeights_4_1 = io_inConf_bits_confneuralNetsinputWeights_4_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_inputWeights_4_2 = io_inConf_bits_confneuralNetsinputWeights_4_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_inputWeights_4_3 = io_inConf_bits_confneuralNetsinputWeights_4_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_inputWeights_5_0 = io_inConf_bits_confneuralNetsinputWeights_5_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_inputWeights_5_1 = io_inConf_bits_confneuralNetsinputWeights_5_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_inputWeights_5_2 = io_inConf_bits_confneuralNetsinputWeights_5_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_inputWeights_5_3 = io_inConf_bits_confneuralNetsinputWeights_5_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_inputWeights_6_0 = io_inConf_bits_confneuralNetsinputWeights_6_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_inputWeights_6_1 = io_inConf_bits_confneuralNetsinputWeights_6_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_inputWeights_6_2 = io_inConf_bits_confneuralNetsinputWeights_6_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_inputWeights_6_3 = io_inConf_bits_confneuralNetsinputWeights_6_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_inputWeights_7_0 = io_inConf_bits_confneuralNetsinputWeights_7_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_inputWeights_7_1 = io_inConf_bits_confneuralNetsinputWeights_7_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_inputWeights_7_2 = io_inConf_bits_confneuralNetsinputWeights_7_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_inputWeights_7_3 = io_inConf_bits_confneuralNetsinputWeights_7_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_inputWeights_8_0 = io_inConf_bits_confneuralNetsinputWeights_8_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_inputWeights_8_1 = io_inConf_bits_confneuralNetsinputWeights_8_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_inputWeights_8_2 = io_inConf_bits_confneuralNetsinputWeights_8_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_inputWeights_8_3 = io_inConf_bits_confneuralNetsinputWeights_8_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_inputWeights_9_0 = io_inConf_bits_confneuralNetsinputWeights_9_0; // @[Wellness.scala 336:30]
  assign neuralNets_io_inputWeights_9_1 = io_inConf_bits_confneuralNetsinputWeights_9_1; // @[Wellness.scala 336:30]
  assign neuralNets_io_inputWeights_9_2 = io_inConf_bits_confneuralNetsinputWeights_9_2; // @[Wellness.scala 336:30]
  assign neuralNets_io_inputWeights_9_3 = io_inConf_bits_confneuralNetsinputWeights_9_3; // @[Wellness.scala 336:30]
  assign neuralNets_io_midAndOutputWeights_0_0 = io_inConf_bits_confneuralNetsmidAndOutputWeights_0_0; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_0_1 = io_inConf_bits_confneuralNetsmidAndOutputWeights_0_1; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_0_2 = io_inConf_bits_confneuralNetsmidAndOutputWeights_0_2; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_0_3 = io_inConf_bits_confneuralNetsmidAndOutputWeights_0_3; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_0_4 = io_inConf_bits_confneuralNetsmidAndOutputWeights_0_4; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_0_5 = io_inConf_bits_confneuralNetsmidAndOutputWeights_0_5; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_0_6 = io_inConf_bits_confneuralNetsmidAndOutputWeights_0_6; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_0_7 = io_inConf_bits_confneuralNetsmidAndOutputWeights_0_7; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_0_8 = io_inConf_bits_confneuralNetsmidAndOutputWeights_0_8; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_0_9 = io_inConf_bits_confneuralNetsmidAndOutputWeights_0_9; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_1_0 = io_inConf_bits_confneuralNetsmidAndOutputWeights_1_0; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_1_1 = io_inConf_bits_confneuralNetsmidAndOutputWeights_1_1; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_1_2 = io_inConf_bits_confneuralNetsmidAndOutputWeights_1_2; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_1_3 = io_inConf_bits_confneuralNetsmidAndOutputWeights_1_3; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_1_4 = io_inConf_bits_confneuralNetsmidAndOutputWeights_1_4; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_1_5 = io_inConf_bits_confneuralNetsmidAndOutputWeights_1_5; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_1_6 = io_inConf_bits_confneuralNetsmidAndOutputWeights_1_6; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_1_7 = io_inConf_bits_confneuralNetsmidAndOutputWeights_1_7; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_1_8 = io_inConf_bits_confneuralNetsmidAndOutputWeights_1_8; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_1_9 = io_inConf_bits_confneuralNetsmidAndOutputWeights_1_9; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_2_0 = io_inConf_bits_confneuralNetsmidAndOutputWeights_2_0; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_2_1 = io_inConf_bits_confneuralNetsmidAndOutputWeights_2_1; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_2_2 = io_inConf_bits_confneuralNetsmidAndOutputWeights_2_2; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_2_3 = io_inConf_bits_confneuralNetsmidAndOutputWeights_2_3; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_2_4 = io_inConf_bits_confneuralNetsmidAndOutputWeights_2_4; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_2_5 = io_inConf_bits_confneuralNetsmidAndOutputWeights_2_5; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_2_6 = io_inConf_bits_confneuralNetsmidAndOutputWeights_2_6; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_2_7 = io_inConf_bits_confneuralNetsmidAndOutputWeights_2_7; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_2_8 = io_inConf_bits_confneuralNetsmidAndOutputWeights_2_8; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_2_9 = io_inConf_bits_confneuralNetsmidAndOutputWeights_2_9; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_3_0 = io_inConf_bits_confneuralNetsmidAndOutputWeights_3_0; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_3_1 = io_inConf_bits_confneuralNetsmidAndOutputWeights_3_1; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_3_2 = io_inConf_bits_confneuralNetsmidAndOutputWeights_3_2; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_3_3 = io_inConf_bits_confneuralNetsmidAndOutputWeights_3_3; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_3_4 = io_inConf_bits_confneuralNetsmidAndOutputWeights_3_4; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_3_5 = io_inConf_bits_confneuralNetsmidAndOutputWeights_3_5; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_3_6 = io_inConf_bits_confneuralNetsmidAndOutputWeights_3_6; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_3_7 = io_inConf_bits_confneuralNetsmidAndOutputWeights_3_7; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_3_8 = io_inConf_bits_confneuralNetsmidAndOutputWeights_3_8; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_3_9 = io_inConf_bits_confneuralNetsmidAndOutputWeights_3_9; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_4_0 = io_inConf_bits_confneuralNetsmidAndOutputWeights_4_0; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_4_1 = io_inConf_bits_confneuralNetsmidAndOutputWeights_4_1; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_4_2 = io_inConf_bits_confneuralNetsmidAndOutputWeights_4_2; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_4_3 = io_inConf_bits_confneuralNetsmidAndOutputWeights_4_3; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_4_4 = io_inConf_bits_confneuralNetsmidAndOutputWeights_4_4; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_4_5 = io_inConf_bits_confneuralNetsmidAndOutputWeights_4_5; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_4_6 = io_inConf_bits_confneuralNetsmidAndOutputWeights_4_6; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_4_7 = io_inConf_bits_confneuralNetsmidAndOutputWeights_4_7; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_4_8 = io_inConf_bits_confneuralNetsmidAndOutputWeights_4_8; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_4_9 = io_inConf_bits_confneuralNetsmidAndOutputWeights_4_9; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_5_0 = io_inConf_bits_confneuralNetsmidAndOutputWeights_5_0; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_5_1 = io_inConf_bits_confneuralNetsmidAndOutputWeights_5_1; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_5_2 = io_inConf_bits_confneuralNetsmidAndOutputWeights_5_2; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_5_3 = io_inConf_bits_confneuralNetsmidAndOutputWeights_5_3; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_5_4 = io_inConf_bits_confneuralNetsmidAndOutputWeights_5_4; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_5_5 = io_inConf_bits_confneuralNetsmidAndOutputWeights_5_5; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_5_6 = io_inConf_bits_confneuralNetsmidAndOutputWeights_5_6; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_5_7 = io_inConf_bits_confneuralNetsmidAndOutputWeights_5_7; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_5_8 = io_inConf_bits_confneuralNetsmidAndOutputWeights_5_8; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_5_9 = io_inConf_bits_confneuralNetsmidAndOutputWeights_5_9; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_6_0 = io_inConf_bits_confneuralNetsmidAndOutputWeights_6_0; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_6_1 = io_inConf_bits_confneuralNetsmidAndOutputWeights_6_1; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_6_2 = io_inConf_bits_confneuralNetsmidAndOutputWeights_6_2; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_6_3 = io_inConf_bits_confneuralNetsmidAndOutputWeights_6_3; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_6_4 = io_inConf_bits_confneuralNetsmidAndOutputWeights_6_4; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_6_5 = io_inConf_bits_confneuralNetsmidAndOutputWeights_6_5; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_6_6 = io_inConf_bits_confneuralNetsmidAndOutputWeights_6_6; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_6_7 = io_inConf_bits_confneuralNetsmidAndOutputWeights_6_7; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_6_8 = io_inConf_bits_confneuralNetsmidAndOutputWeights_6_8; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_6_9 = io_inConf_bits_confneuralNetsmidAndOutputWeights_6_9; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_7_0 = io_inConf_bits_confneuralNetsmidAndOutputWeights_7_0; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_7_1 = io_inConf_bits_confneuralNetsmidAndOutputWeights_7_1; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_7_2 = io_inConf_bits_confneuralNetsmidAndOutputWeights_7_2; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_7_3 = io_inConf_bits_confneuralNetsmidAndOutputWeights_7_3; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_7_4 = io_inConf_bits_confneuralNetsmidAndOutputWeights_7_4; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_7_5 = io_inConf_bits_confneuralNetsmidAndOutputWeights_7_5; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_7_6 = io_inConf_bits_confneuralNetsmidAndOutputWeights_7_6; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_7_7 = io_inConf_bits_confneuralNetsmidAndOutputWeights_7_7; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_7_8 = io_inConf_bits_confneuralNetsmidAndOutputWeights_7_8; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_7_9 = io_inConf_bits_confneuralNetsmidAndOutputWeights_7_9; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_8_0 = io_inConf_bits_confneuralNetsmidAndOutputWeights_8_0; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_8_1 = io_inConf_bits_confneuralNetsmidAndOutputWeights_8_1; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_8_2 = io_inConf_bits_confneuralNetsmidAndOutputWeights_8_2; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_8_3 = io_inConf_bits_confneuralNetsmidAndOutputWeights_8_3; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_8_4 = io_inConf_bits_confneuralNetsmidAndOutputWeights_8_4; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_8_5 = io_inConf_bits_confneuralNetsmidAndOutputWeights_8_5; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_8_6 = io_inConf_bits_confneuralNetsmidAndOutputWeights_8_6; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_8_7 = io_inConf_bits_confneuralNetsmidAndOutputWeights_8_7; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_8_8 = io_inConf_bits_confneuralNetsmidAndOutputWeights_8_8; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_8_9 = io_inConf_bits_confneuralNetsmidAndOutputWeights_8_9; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_9_0 = io_inConf_bits_confneuralNetsmidAndOutputWeights_9_0; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_9_1 = io_inConf_bits_confneuralNetsmidAndOutputWeights_9_1; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_9_2 = io_inConf_bits_confneuralNetsmidAndOutputWeights_9_2; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_9_3 = io_inConf_bits_confneuralNetsmidAndOutputWeights_9_3; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_9_4 = io_inConf_bits_confneuralNetsmidAndOutputWeights_9_4; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_9_5 = io_inConf_bits_confneuralNetsmidAndOutputWeights_9_5; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_9_6 = io_inConf_bits_confneuralNetsmidAndOutputWeights_9_6; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_9_7 = io_inConf_bits_confneuralNetsmidAndOutputWeights_9_7; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_9_8 = io_inConf_bits_confneuralNetsmidAndOutputWeights_9_8; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_9_9 = io_inConf_bits_confneuralNetsmidAndOutputWeights_9_9; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_10_0 = io_inConf_bits_confneuralNetsmidAndOutputWeights_10_0; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_10_1 = io_inConf_bits_confneuralNetsmidAndOutputWeights_10_1; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_10_2 = io_inConf_bits_confneuralNetsmidAndOutputWeights_10_2; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_10_3 = io_inConf_bits_confneuralNetsmidAndOutputWeights_10_3; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_10_4 = io_inConf_bits_confneuralNetsmidAndOutputWeights_10_4; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_10_5 = io_inConf_bits_confneuralNetsmidAndOutputWeights_10_5; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_10_6 = io_inConf_bits_confneuralNetsmidAndOutputWeights_10_6; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_10_7 = io_inConf_bits_confneuralNetsmidAndOutputWeights_10_7; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_10_8 = io_inConf_bits_confneuralNetsmidAndOutputWeights_10_8; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_10_9 = io_inConf_bits_confneuralNetsmidAndOutputWeights_10_9; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_11_0 = io_inConf_bits_confneuralNetsmidAndOutputWeights_11_0; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_11_1 = io_inConf_bits_confneuralNetsmidAndOutputWeights_11_1; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_11_2 = io_inConf_bits_confneuralNetsmidAndOutputWeights_11_2; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_11_3 = io_inConf_bits_confneuralNetsmidAndOutputWeights_11_3; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_11_4 = io_inConf_bits_confneuralNetsmidAndOutputWeights_11_4; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_11_5 = io_inConf_bits_confneuralNetsmidAndOutputWeights_11_5; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_11_6 = io_inConf_bits_confneuralNetsmidAndOutputWeights_11_6; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_11_7 = io_inConf_bits_confneuralNetsmidAndOutputWeights_11_7; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_11_8 = io_inConf_bits_confneuralNetsmidAndOutputWeights_11_8; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_11_9 = io_inConf_bits_confneuralNetsmidAndOutputWeights_11_9; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_12_0 = io_inConf_bits_confneuralNetsmidAndOutputWeights_12_0; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_12_1 = io_inConf_bits_confneuralNetsmidAndOutputWeights_12_1; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_12_2 = io_inConf_bits_confneuralNetsmidAndOutputWeights_12_2; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_12_3 = io_inConf_bits_confneuralNetsmidAndOutputWeights_12_3; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_12_4 = io_inConf_bits_confneuralNetsmidAndOutputWeights_12_4; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_12_5 = io_inConf_bits_confneuralNetsmidAndOutputWeights_12_5; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_12_6 = io_inConf_bits_confneuralNetsmidAndOutputWeights_12_6; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_12_7 = io_inConf_bits_confneuralNetsmidAndOutputWeights_12_7; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_12_8 = io_inConf_bits_confneuralNetsmidAndOutputWeights_12_8; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_12_9 = io_inConf_bits_confneuralNetsmidAndOutputWeights_12_9; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_13_0 = io_inConf_bits_confneuralNetsmidAndOutputWeights_13_0; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_13_1 = io_inConf_bits_confneuralNetsmidAndOutputWeights_13_1; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_13_2 = io_inConf_bits_confneuralNetsmidAndOutputWeights_13_2; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_13_3 = io_inConf_bits_confneuralNetsmidAndOutputWeights_13_3; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_13_4 = io_inConf_bits_confneuralNetsmidAndOutputWeights_13_4; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_13_5 = io_inConf_bits_confneuralNetsmidAndOutputWeights_13_5; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_13_6 = io_inConf_bits_confneuralNetsmidAndOutputWeights_13_6; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_13_7 = io_inConf_bits_confneuralNetsmidAndOutputWeights_13_7; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_13_8 = io_inConf_bits_confneuralNetsmidAndOutputWeights_13_8; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_13_9 = io_inConf_bits_confneuralNetsmidAndOutputWeights_13_9; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_14_0 = io_inConf_bits_confneuralNetsmidAndOutputWeights_14_0; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_14_1 = io_inConf_bits_confneuralNetsmidAndOutputWeights_14_1; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_14_2 = io_inConf_bits_confneuralNetsmidAndOutputWeights_14_2; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_14_3 = io_inConf_bits_confneuralNetsmidAndOutputWeights_14_3; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_14_4 = io_inConf_bits_confneuralNetsmidAndOutputWeights_14_4; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_14_5 = io_inConf_bits_confneuralNetsmidAndOutputWeights_14_5; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_14_6 = io_inConf_bits_confneuralNetsmidAndOutputWeights_14_6; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_14_7 = io_inConf_bits_confneuralNetsmidAndOutputWeights_14_7; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_14_8 = io_inConf_bits_confneuralNetsmidAndOutputWeights_14_8; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_14_9 = io_inConf_bits_confneuralNetsmidAndOutputWeights_14_9; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_15_0 = io_inConf_bits_confneuralNetsmidAndOutputWeights_15_0; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_15_1 = io_inConf_bits_confneuralNetsmidAndOutputWeights_15_1; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_15_2 = io_inConf_bits_confneuralNetsmidAndOutputWeights_15_2; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_15_3 = io_inConf_bits_confneuralNetsmidAndOutputWeights_15_3; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_15_4 = io_inConf_bits_confneuralNetsmidAndOutputWeights_15_4; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_15_5 = io_inConf_bits_confneuralNetsmidAndOutputWeights_15_5; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_15_6 = io_inConf_bits_confneuralNetsmidAndOutputWeights_15_6; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_15_7 = io_inConf_bits_confneuralNetsmidAndOutputWeights_15_7; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_15_8 = io_inConf_bits_confneuralNetsmidAndOutputWeights_15_8; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_15_9 = io_inConf_bits_confneuralNetsmidAndOutputWeights_15_9; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_16_0 = io_inConf_bits_confneuralNetsmidAndOutputWeights_16_0; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_16_1 = io_inConf_bits_confneuralNetsmidAndOutputWeights_16_1; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_16_2 = io_inConf_bits_confneuralNetsmidAndOutputWeights_16_2; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_16_3 = io_inConf_bits_confneuralNetsmidAndOutputWeights_16_3; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_16_4 = io_inConf_bits_confneuralNetsmidAndOutputWeights_16_4; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_16_5 = io_inConf_bits_confneuralNetsmidAndOutputWeights_16_5; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_16_6 = io_inConf_bits_confneuralNetsmidAndOutputWeights_16_6; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_16_7 = io_inConf_bits_confneuralNetsmidAndOutputWeights_16_7; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_16_8 = io_inConf_bits_confneuralNetsmidAndOutputWeights_16_8; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_16_9 = io_inConf_bits_confneuralNetsmidAndOutputWeights_16_9; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_17_0 = io_inConf_bits_confneuralNetsmidAndOutputWeights_17_0; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_17_1 = io_inConf_bits_confneuralNetsmidAndOutputWeights_17_1; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_17_2 = io_inConf_bits_confneuralNetsmidAndOutputWeights_17_2; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_17_3 = io_inConf_bits_confneuralNetsmidAndOutputWeights_17_3; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_17_4 = io_inConf_bits_confneuralNetsmidAndOutputWeights_17_4; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_17_5 = io_inConf_bits_confneuralNetsmidAndOutputWeights_17_5; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_17_6 = io_inConf_bits_confneuralNetsmidAndOutputWeights_17_6; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_17_7 = io_inConf_bits_confneuralNetsmidAndOutputWeights_17_7; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_17_8 = io_inConf_bits_confneuralNetsmidAndOutputWeights_17_8; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_17_9 = io_inConf_bits_confneuralNetsmidAndOutputWeights_17_9; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_18_0 = io_inConf_bits_confneuralNetsmidAndOutputWeights_18_0; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_18_1 = io_inConf_bits_confneuralNetsmidAndOutputWeights_18_1; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_18_2 = io_inConf_bits_confneuralNetsmidAndOutputWeights_18_2; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_18_3 = io_inConf_bits_confneuralNetsmidAndOutputWeights_18_3; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_18_4 = io_inConf_bits_confneuralNetsmidAndOutputWeights_18_4; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_18_5 = io_inConf_bits_confneuralNetsmidAndOutputWeights_18_5; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_18_6 = io_inConf_bits_confneuralNetsmidAndOutputWeights_18_6; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_18_7 = io_inConf_bits_confneuralNetsmidAndOutputWeights_18_7; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_18_8 = io_inConf_bits_confneuralNetsmidAndOutputWeights_18_8; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_18_9 = io_inConf_bits_confneuralNetsmidAndOutputWeights_18_9; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_19_0 = io_inConf_bits_confneuralNetsmidAndOutputWeights_19_0; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_19_1 = io_inConf_bits_confneuralNetsmidAndOutputWeights_19_1; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_19_2 = io_inConf_bits_confneuralNetsmidAndOutputWeights_19_2; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_19_3 = io_inConf_bits_confneuralNetsmidAndOutputWeights_19_3; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_19_4 = io_inConf_bits_confneuralNetsmidAndOutputWeights_19_4; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_19_5 = io_inConf_bits_confneuralNetsmidAndOutputWeights_19_5; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_19_6 = io_inConf_bits_confneuralNetsmidAndOutputWeights_19_6; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_19_7 = io_inConf_bits_confneuralNetsmidAndOutputWeights_19_7; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_19_8 = io_inConf_bits_confneuralNetsmidAndOutputWeights_19_8; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_19_9 = io_inConf_bits_confneuralNetsmidAndOutputWeights_19_9; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_20_0 = io_inConf_bits_confneuralNetsmidAndOutputWeights_20_0; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_20_1 = io_inConf_bits_confneuralNetsmidAndOutputWeights_20_1; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_20_2 = io_inConf_bits_confneuralNetsmidAndOutputWeights_20_2; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_20_3 = io_inConf_bits_confneuralNetsmidAndOutputWeights_20_3; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_20_4 = io_inConf_bits_confneuralNetsmidAndOutputWeights_20_4; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_20_5 = io_inConf_bits_confneuralNetsmidAndOutputWeights_20_5; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_20_6 = io_inConf_bits_confneuralNetsmidAndOutputWeights_20_6; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_20_7 = io_inConf_bits_confneuralNetsmidAndOutputWeights_20_7; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_20_8 = io_inConf_bits_confneuralNetsmidAndOutputWeights_20_8; // @[Wellness.scala 337:37]
  assign neuralNets_io_midAndOutputWeights_20_9 = io_inConf_bits_confneuralNetsmidAndOutputWeights_20_9; // @[Wellness.scala 337:37]
  assign neuralNets_io_biasVecs_0_0 = io_inConf_bits_confneuralNetsbiasVecs_0_0; // @[Wellness.scala 338:26]
  assign neuralNets_io_biasVecs_0_1 = io_inConf_bits_confneuralNetsbiasVecs_0_1; // @[Wellness.scala 338:26]
  assign neuralNets_io_biasVecs_0_2 = io_inConf_bits_confneuralNetsbiasVecs_0_2; // @[Wellness.scala 338:26]
  assign neuralNets_io_biasVecs_0_3 = io_inConf_bits_confneuralNetsbiasVecs_0_3; // @[Wellness.scala 338:26]
  assign neuralNets_io_biasVecs_0_4 = io_inConf_bits_confneuralNetsbiasVecs_0_4; // @[Wellness.scala 338:26]
  assign neuralNets_io_biasVecs_0_5 = io_inConf_bits_confneuralNetsbiasVecs_0_5; // @[Wellness.scala 338:26]
  assign neuralNets_io_biasVecs_0_6 = io_inConf_bits_confneuralNetsbiasVecs_0_6; // @[Wellness.scala 338:26]
  assign neuralNets_io_biasVecs_0_7 = io_inConf_bits_confneuralNetsbiasVecs_0_7; // @[Wellness.scala 338:26]
  assign neuralNets_io_biasVecs_0_8 = io_inConf_bits_confneuralNetsbiasVecs_0_8; // @[Wellness.scala 338:26]
  assign neuralNets_io_biasVecs_0_9 = io_inConf_bits_confneuralNetsbiasVecs_0_9; // @[Wellness.scala 338:26]
  assign neuralNets_io_biasVecs_1_0 = io_inConf_bits_confneuralNetsbiasVecs_1_0; // @[Wellness.scala 338:26]
  assign neuralNets_io_biasVecs_1_1 = io_inConf_bits_confneuralNetsbiasVecs_1_1; // @[Wellness.scala 338:26]
  assign neuralNets_io_biasVecs_1_2 = io_inConf_bits_confneuralNetsbiasVecs_1_2; // @[Wellness.scala 338:26]
  assign neuralNets_io_biasVecs_1_3 = io_inConf_bits_confneuralNetsbiasVecs_1_3; // @[Wellness.scala 338:26]
  assign neuralNets_io_biasVecs_1_4 = io_inConf_bits_confneuralNetsbiasVecs_1_4; // @[Wellness.scala 338:26]
  assign neuralNets_io_biasVecs_1_5 = io_inConf_bits_confneuralNetsbiasVecs_1_5; // @[Wellness.scala 338:26]
  assign neuralNets_io_biasVecs_1_6 = io_inConf_bits_confneuralNetsbiasVecs_1_6; // @[Wellness.scala 338:26]
  assign neuralNets_io_biasVecs_1_7 = io_inConf_bits_confneuralNetsbiasVecs_1_7; // @[Wellness.scala 338:26]
  assign neuralNets_io_biasVecs_1_8 = io_inConf_bits_confneuralNetsbiasVecs_1_8; // @[Wellness.scala 338:26]
  assign neuralNets_io_biasVecs_1_9 = io_inConf_bits_confneuralNetsbiasVecs_1_9; // @[Wellness.scala 338:26]
  assign neuralNets_io_biasVecs_2_0 = io_inConf_bits_confneuralNetsbiasVecs_2_0; // @[Wellness.scala 338:26]
  assign neuralNets_io_biasVecs_2_1 = io_inConf_bits_confneuralNetsbiasVecs_2_1; // @[Wellness.scala 338:26]
  assign neuralNets_io_biasVecs_2_2 = io_inConf_bits_confneuralNetsbiasVecs_2_2; // @[Wellness.scala 338:26]
  assign neuralNets_io_biasVecs_2_3 = io_inConf_bits_confneuralNetsbiasVecs_2_3; // @[Wellness.scala 338:26]
  assign neuralNets_io_biasVecs_2_4 = io_inConf_bits_confneuralNetsbiasVecs_2_4; // @[Wellness.scala 338:26]
  assign neuralNets_io_biasVecs_2_5 = io_inConf_bits_confneuralNetsbiasVecs_2_5; // @[Wellness.scala 338:26]
  assign neuralNets_io_biasVecs_2_6 = io_inConf_bits_confneuralNetsbiasVecs_2_6; // @[Wellness.scala 338:26]
  assign neuralNets_io_biasVecs_2_7 = io_inConf_bits_confneuralNetsbiasVecs_2_7; // @[Wellness.scala 338:26]
  assign neuralNets_io_biasVecs_2_8 = io_inConf_bits_confneuralNetsbiasVecs_2_8; // @[Wellness.scala 338:26]
  assign neuralNets_io_biasVecs_2_9 = io_inConf_bits_confneuralNetsbiasVecs_2_9; // @[Wellness.scala 338:26]
  assign neuralNets_io_outputBias = io_inConf_bits_confneuralNetsoutputBias_0; // @[Wellness.scala 339:28]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  lineLength1Reg1 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  lineLength1Valid1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    lineLength1Reg1 <= $signed(_T_22);
    lineLength1Valid1 <= lineLength1_io_out_valid;
  end
endmodule
module MemoryBuffer(
  input         clock,
  input         reset,
  input         io_in_valid,
  input  [31:0] io_in_bits,
  output [31:0] io_out_bits_0_0,
  output [31:0] io_out_bits_0_1,
  output [31:0] io_out_bits_0_2,
  output [31:0] io_out_bits_0_3,
  output [31:0] io_out_bits_1_0,
  output [31:0] io_out_bits_1_1,
  output [31:0] io_out_bits_1_2,
  output [31:0] io_out_bits_1_3,
  output [31:0] io_out_bits_2_0,
  output [31:0] io_out_bits_2_1,
  output [31:0] io_out_bits_2_2,
  output [31:0] io_out_bits_2_3,
  output [31:0] io_out_bits_3_0,
  output [31:0] io_out_bits_3_1,
  output [31:0] io_out_bits_3_2,
  output [31:0] io_out_bits_3_3,
  output [31:0] io_out_bits_4_0,
  output [31:0] io_out_bits_4_1,
  output [31:0] io_out_bits_4_2,
  output [31:0] io_out_bits_4_3,
  output [31:0] io_out_bits_5_0,
  output [31:0] io_out_bits_5_1,
  output [31:0] io_out_bits_5_2,
  output [31:0] io_out_bits_5_3,
  output [31:0] io_out_bits_6_0,
  output [31:0] io_out_bits_6_1,
  output [31:0] io_out_bits_6_2,
  output [31:0] io_out_bits_6_3,
  output [31:0] io_out_bits_7_0,
  output [31:0] io_out_bits_7_1,
  output [31:0] io_out_bits_7_2,
  output [31:0] io_out_bits_7_3,
  output [31:0] io_out_bits_8_0,
  output [31:0] io_out_bits_8_1,
  output [31:0] io_out_bits_8_2,
  output [31:0] io_out_bits_8_3,
  output [31:0] io_out_bits_9_0,
  output [31:0] io_out_bits_9_1,
  output [31:0] io_out_bits_9_2,
  output [31:0] io_out_bits_9_3
);
  reg [31:0] regs_0; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_0;
  reg [31:0] regs_1; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_1;
  reg [31:0] regs_2; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_2;
  reg [31:0] regs_3; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_3;
  reg [31:0] regs_4; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_4;
  reg [31:0] regs_5; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_5;
  reg [31:0] regs_6; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_6;
  reg [31:0] regs_7; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_7;
  reg [31:0] regs_8; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_8;
  reg [31:0] regs_9; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_9;
  reg [31:0] regs_10; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_10;
  reg [31:0] regs_11; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_11;
  reg [31:0] regs_12; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_12;
  reg [31:0] regs_13; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_13;
  reg [31:0] regs_14; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_14;
  reg [31:0] regs_15; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_15;
  reg [31:0] regs_16; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_16;
  reg [31:0] regs_17; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_17;
  reg [31:0] regs_18; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_18;
  reg [31:0] regs_19; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_19;
  reg [31:0] regs_20; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_20;
  reg [31:0] regs_21; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_21;
  reg [31:0] regs_22; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_22;
  reg [31:0] regs_23; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_23;
  reg [31:0] regs_24; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_24;
  reg [31:0] regs_25; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_25;
  reg [31:0] regs_26; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_26;
  reg [31:0] regs_27; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_27;
  reg [31:0] regs_28; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_28;
  reg [31:0] regs_29; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_29;
  reg [31:0] regs_30; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_30;
  reg [31:0] regs_31; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_31;
  reg [31:0] regs_32; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_32;
  reg [31:0] regs_33; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_33;
  reg [31:0] regs_34; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_34;
  reg [31:0] regs_35; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_35;
  reg [31:0] regs_36; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_36;
  reg [31:0] regs_37; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_37;
  reg [31:0] regs_38; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_38;
  reg [31:0] regs_39; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_39;
  assign io_out_bits_0_0 = regs_0; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_1 = regs_1; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_2 = regs_2; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_3 = regs_3; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_1_0 = regs_4; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_1_1 = regs_5; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_1_2 = regs_6; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_1_3 = regs_7; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_2_0 = regs_8; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_2_1 = regs_9; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_2_2 = regs_10; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_2_3 = regs_11; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_3_0 = regs_12; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_3_1 = regs_13; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_3_2 = regs_14; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_3_3 = regs_15; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_4_0 = regs_16; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_4_1 = regs_17; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_4_2 = regs_18; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_4_3 = regs_19; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_5_0 = regs_20; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_5_1 = regs_21; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_5_2 = regs_22; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_5_3 = regs_23; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_6_0 = regs_24; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_6_1 = regs_25; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_6_2 = regs_26; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_6_3 = regs_27; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_7_0 = regs_28; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_7_1 = regs_29; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_7_2 = regs_30; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_7_3 = regs_31; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_8_0 = regs_32; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_8_1 = regs_33; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_8_2 = regs_34; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_8_3 = regs_35; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_9_0 = regs_36; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_9_1 = regs_37; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_9_2 = regs_38; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_9_3 = regs_39; // @[MemoryBuffer.scala 65:25]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  regs_3 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  regs_4 = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  regs_5 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  regs_6 = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  regs_7 = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  regs_8 = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  regs_9 = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  regs_10 = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  regs_11 = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  regs_12 = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  regs_13 = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  regs_14 = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  regs_15 = _RAND_15[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  regs_16 = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  regs_17 = _RAND_17[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  regs_18 = _RAND_18[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  regs_19 = _RAND_19[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  regs_20 = _RAND_20[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  regs_21 = _RAND_21[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  regs_22 = _RAND_22[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  regs_23 = _RAND_23[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  regs_24 = _RAND_24[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  regs_25 = _RAND_25[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  regs_26 = _RAND_26[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  regs_27 = _RAND_27[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  regs_28 = _RAND_28[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  regs_29 = _RAND_29[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  regs_30 = _RAND_30[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  regs_31 = _RAND_31[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  regs_32 = _RAND_32[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  regs_33 = _RAND_33[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  regs_34 = _RAND_34[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  regs_35 = _RAND_35[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  regs_36 = _RAND_36[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  regs_37 = _RAND_37[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  regs_38 = _RAND_38[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  regs_39 = _RAND_39[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      regs_0 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_0 <= io_in_bits;
      end
    end
    if (reset) begin
      regs_1 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_1 <= regs_0;
      end
    end
    if (reset) begin
      regs_2 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_2 <= regs_1;
      end
    end
    if (reset) begin
      regs_3 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_3 <= regs_2;
      end
    end
    if (reset) begin
      regs_4 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_4 <= regs_3;
      end
    end
    if (reset) begin
      regs_5 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_5 <= regs_4;
      end
    end
    if (reset) begin
      regs_6 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_6 <= regs_5;
      end
    end
    if (reset) begin
      regs_7 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_7 <= regs_6;
      end
    end
    if (reset) begin
      regs_8 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_8 <= regs_7;
      end
    end
    if (reset) begin
      regs_9 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_9 <= regs_8;
      end
    end
    if (reset) begin
      regs_10 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_10 <= regs_9;
      end
    end
    if (reset) begin
      regs_11 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_11 <= regs_10;
      end
    end
    if (reset) begin
      regs_12 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_12 <= regs_11;
      end
    end
    if (reset) begin
      regs_13 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_13 <= regs_12;
      end
    end
    if (reset) begin
      regs_14 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_14 <= regs_13;
      end
    end
    if (reset) begin
      regs_15 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_15 <= regs_14;
      end
    end
    if (reset) begin
      regs_16 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_16 <= regs_15;
      end
    end
    if (reset) begin
      regs_17 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_17 <= regs_16;
      end
    end
    if (reset) begin
      regs_18 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_18 <= regs_17;
      end
    end
    if (reset) begin
      regs_19 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_19 <= regs_18;
      end
    end
    if (reset) begin
      regs_20 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_20 <= regs_19;
      end
    end
    if (reset) begin
      regs_21 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_21 <= regs_20;
      end
    end
    if (reset) begin
      regs_22 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_22 <= regs_21;
      end
    end
    if (reset) begin
      regs_23 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_23 <= regs_22;
      end
    end
    if (reset) begin
      regs_24 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_24 <= regs_23;
      end
    end
    if (reset) begin
      regs_25 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_25 <= regs_24;
      end
    end
    if (reset) begin
      regs_26 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_26 <= regs_25;
      end
    end
    if (reset) begin
      regs_27 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_27 <= regs_26;
      end
    end
    if (reset) begin
      regs_28 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_28 <= regs_27;
      end
    end
    if (reset) begin
      regs_29 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_29 <= regs_28;
      end
    end
    if (reset) begin
      regs_30 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_30 <= regs_29;
      end
    end
    if (reset) begin
      regs_31 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_31 <= regs_30;
      end
    end
    if (reset) begin
      regs_32 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_32 <= regs_31;
      end
    end
    if (reset) begin
      regs_33 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_33 <= regs_32;
      end
    end
    if (reset) begin
      regs_34 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_34 <= regs_33;
      end
    end
    if (reset) begin
      regs_35 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_35 <= regs_34;
      end
    end
    if (reset) begin
      regs_36 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_36 <= regs_35;
      end
    end
    if (reset) begin
      regs_37 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_37 <= regs_36;
      end
    end
    if (reset) begin
      regs_38 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_38 <= regs_37;
      end
    end
    if (reset) begin
      regs_39 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_39 <= regs_38;
      end
    end
  end
endmodule
module MemoryBuffer_1(
  input         clock,
  input         reset,
  input         io_in_valid,
  input  [31:0] io_in_bits,
  output [31:0] io_out_bits_0_0,
  output [31:0] io_out_bits_0_1,
  output [31:0] io_out_bits_0_2,
  output [31:0] io_out_bits_0_3,
  output [31:0] io_out_bits_0_4,
  output [31:0] io_out_bits_0_5,
  output [31:0] io_out_bits_0_6,
  output [31:0] io_out_bits_0_7,
  output [31:0] io_out_bits_0_8,
  output [31:0] io_out_bits_0_9,
  output [31:0] io_out_bits_1_0,
  output [31:0] io_out_bits_1_1,
  output [31:0] io_out_bits_1_2,
  output [31:0] io_out_bits_1_3,
  output [31:0] io_out_bits_1_4,
  output [31:0] io_out_bits_1_5,
  output [31:0] io_out_bits_1_6,
  output [31:0] io_out_bits_1_7,
  output [31:0] io_out_bits_1_8,
  output [31:0] io_out_bits_1_9,
  output [31:0] io_out_bits_2_0,
  output [31:0] io_out_bits_2_1,
  output [31:0] io_out_bits_2_2,
  output [31:0] io_out_bits_2_3,
  output [31:0] io_out_bits_2_4,
  output [31:0] io_out_bits_2_5,
  output [31:0] io_out_bits_2_6,
  output [31:0] io_out_bits_2_7,
  output [31:0] io_out_bits_2_8,
  output [31:0] io_out_bits_2_9,
  output [31:0] io_out_bits_3_0,
  output [31:0] io_out_bits_3_1,
  output [31:0] io_out_bits_3_2,
  output [31:0] io_out_bits_3_3,
  output [31:0] io_out_bits_3_4,
  output [31:0] io_out_bits_3_5,
  output [31:0] io_out_bits_3_6,
  output [31:0] io_out_bits_3_7,
  output [31:0] io_out_bits_3_8,
  output [31:0] io_out_bits_3_9,
  output [31:0] io_out_bits_4_0,
  output [31:0] io_out_bits_4_1,
  output [31:0] io_out_bits_4_2,
  output [31:0] io_out_bits_4_3,
  output [31:0] io_out_bits_4_4,
  output [31:0] io_out_bits_4_5,
  output [31:0] io_out_bits_4_6,
  output [31:0] io_out_bits_4_7,
  output [31:0] io_out_bits_4_8,
  output [31:0] io_out_bits_4_9,
  output [31:0] io_out_bits_5_0,
  output [31:0] io_out_bits_5_1,
  output [31:0] io_out_bits_5_2,
  output [31:0] io_out_bits_5_3,
  output [31:0] io_out_bits_5_4,
  output [31:0] io_out_bits_5_5,
  output [31:0] io_out_bits_5_6,
  output [31:0] io_out_bits_5_7,
  output [31:0] io_out_bits_5_8,
  output [31:0] io_out_bits_5_9,
  output [31:0] io_out_bits_6_0,
  output [31:0] io_out_bits_6_1,
  output [31:0] io_out_bits_6_2,
  output [31:0] io_out_bits_6_3,
  output [31:0] io_out_bits_6_4,
  output [31:0] io_out_bits_6_5,
  output [31:0] io_out_bits_6_6,
  output [31:0] io_out_bits_6_7,
  output [31:0] io_out_bits_6_8,
  output [31:0] io_out_bits_6_9,
  output [31:0] io_out_bits_7_0,
  output [31:0] io_out_bits_7_1,
  output [31:0] io_out_bits_7_2,
  output [31:0] io_out_bits_7_3,
  output [31:0] io_out_bits_7_4,
  output [31:0] io_out_bits_7_5,
  output [31:0] io_out_bits_7_6,
  output [31:0] io_out_bits_7_7,
  output [31:0] io_out_bits_7_8,
  output [31:0] io_out_bits_7_9,
  output [31:0] io_out_bits_8_0,
  output [31:0] io_out_bits_8_1,
  output [31:0] io_out_bits_8_2,
  output [31:0] io_out_bits_8_3,
  output [31:0] io_out_bits_8_4,
  output [31:0] io_out_bits_8_5,
  output [31:0] io_out_bits_8_6,
  output [31:0] io_out_bits_8_7,
  output [31:0] io_out_bits_8_8,
  output [31:0] io_out_bits_8_9,
  output [31:0] io_out_bits_9_0,
  output [31:0] io_out_bits_9_1,
  output [31:0] io_out_bits_9_2,
  output [31:0] io_out_bits_9_3,
  output [31:0] io_out_bits_9_4,
  output [31:0] io_out_bits_9_5,
  output [31:0] io_out_bits_9_6,
  output [31:0] io_out_bits_9_7,
  output [31:0] io_out_bits_9_8,
  output [31:0] io_out_bits_9_9,
  output [31:0] io_out_bits_10_0,
  output [31:0] io_out_bits_10_1,
  output [31:0] io_out_bits_10_2,
  output [31:0] io_out_bits_10_3,
  output [31:0] io_out_bits_10_4,
  output [31:0] io_out_bits_10_5,
  output [31:0] io_out_bits_10_6,
  output [31:0] io_out_bits_10_7,
  output [31:0] io_out_bits_10_8,
  output [31:0] io_out_bits_10_9,
  output [31:0] io_out_bits_11_0,
  output [31:0] io_out_bits_11_1,
  output [31:0] io_out_bits_11_2,
  output [31:0] io_out_bits_11_3,
  output [31:0] io_out_bits_11_4,
  output [31:0] io_out_bits_11_5,
  output [31:0] io_out_bits_11_6,
  output [31:0] io_out_bits_11_7,
  output [31:0] io_out_bits_11_8,
  output [31:0] io_out_bits_11_9,
  output [31:0] io_out_bits_12_0,
  output [31:0] io_out_bits_12_1,
  output [31:0] io_out_bits_12_2,
  output [31:0] io_out_bits_12_3,
  output [31:0] io_out_bits_12_4,
  output [31:0] io_out_bits_12_5,
  output [31:0] io_out_bits_12_6,
  output [31:0] io_out_bits_12_7,
  output [31:0] io_out_bits_12_8,
  output [31:0] io_out_bits_12_9,
  output [31:0] io_out_bits_13_0,
  output [31:0] io_out_bits_13_1,
  output [31:0] io_out_bits_13_2,
  output [31:0] io_out_bits_13_3,
  output [31:0] io_out_bits_13_4,
  output [31:0] io_out_bits_13_5,
  output [31:0] io_out_bits_13_6,
  output [31:0] io_out_bits_13_7,
  output [31:0] io_out_bits_13_8,
  output [31:0] io_out_bits_13_9,
  output [31:0] io_out_bits_14_0,
  output [31:0] io_out_bits_14_1,
  output [31:0] io_out_bits_14_2,
  output [31:0] io_out_bits_14_3,
  output [31:0] io_out_bits_14_4,
  output [31:0] io_out_bits_14_5,
  output [31:0] io_out_bits_14_6,
  output [31:0] io_out_bits_14_7,
  output [31:0] io_out_bits_14_8,
  output [31:0] io_out_bits_14_9,
  output [31:0] io_out_bits_15_0,
  output [31:0] io_out_bits_15_1,
  output [31:0] io_out_bits_15_2,
  output [31:0] io_out_bits_15_3,
  output [31:0] io_out_bits_15_4,
  output [31:0] io_out_bits_15_5,
  output [31:0] io_out_bits_15_6,
  output [31:0] io_out_bits_15_7,
  output [31:0] io_out_bits_15_8,
  output [31:0] io_out_bits_15_9,
  output [31:0] io_out_bits_16_0,
  output [31:0] io_out_bits_16_1,
  output [31:0] io_out_bits_16_2,
  output [31:0] io_out_bits_16_3,
  output [31:0] io_out_bits_16_4,
  output [31:0] io_out_bits_16_5,
  output [31:0] io_out_bits_16_6,
  output [31:0] io_out_bits_16_7,
  output [31:0] io_out_bits_16_8,
  output [31:0] io_out_bits_16_9,
  output [31:0] io_out_bits_17_0,
  output [31:0] io_out_bits_17_1,
  output [31:0] io_out_bits_17_2,
  output [31:0] io_out_bits_17_3,
  output [31:0] io_out_bits_17_4,
  output [31:0] io_out_bits_17_5,
  output [31:0] io_out_bits_17_6,
  output [31:0] io_out_bits_17_7,
  output [31:0] io_out_bits_17_8,
  output [31:0] io_out_bits_17_9,
  output [31:0] io_out_bits_18_0,
  output [31:0] io_out_bits_18_1,
  output [31:0] io_out_bits_18_2,
  output [31:0] io_out_bits_18_3,
  output [31:0] io_out_bits_18_4,
  output [31:0] io_out_bits_18_5,
  output [31:0] io_out_bits_18_6,
  output [31:0] io_out_bits_18_7,
  output [31:0] io_out_bits_18_8,
  output [31:0] io_out_bits_18_9,
  output [31:0] io_out_bits_19_0,
  output [31:0] io_out_bits_19_1,
  output [31:0] io_out_bits_19_2,
  output [31:0] io_out_bits_19_3,
  output [31:0] io_out_bits_19_4,
  output [31:0] io_out_bits_19_5,
  output [31:0] io_out_bits_19_6,
  output [31:0] io_out_bits_19_7,
  output [31:0] io_out_bits_19_8,
  output [31:0] io_out_bits_19_9,
  output [31:0] io_out_bits_20_0,
  output [31:0] io_out_bits_20_1,
  output [31:0] io_out_bits_20_2,
  output [31:0] io_out_bits_20_3,
  output [31:0] io_out_bits_20_4,
  output [31:0] io_out_bits_20_5,
  output [31:0] io_out_bits_20_6,
  output [31:0] io_out_bits_20_7,
  output [31:0] io_out_bits_20_8,
  output [31:0] io_out_bits_20_9
);
  reg [31:0] regs_0; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_0;
  reg [31:0] regs_1; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_1;
  reg [31:0] regs_2; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_2;
  reg [31:0] regs_3; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_3;
  reg [31:0] regs_4; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_4;
  reg [31:0] regs_5; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_5;
  reg [31:0] regs_6; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_6;
  reg [31:0] regs_7; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_7;
  reg [31:0] regs_8; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_8;
  reg [31:0] regs_9; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_9;
  reg [31:0] regs_10; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_10;
  reg [31:0] regs_11; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_11;
  reg [31:0] regs_12; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_12;
  reg [31:0] regs_13; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_13;
  reg [31:0] regs_14; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_14;
  reg [31:0] regs_15; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_15;
  reg [31:0] regs_16; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_16;
  reg [31:0] regs_17; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_17;
  reg [31:0] regs_18; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_18;
  reg [31:0] regs_19; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_19;
  reg [31:0] regs_20; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_20;
  reg [31:0] regs_21; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_21;
  reg [31:0] regs_22; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_22;
  reg [31:0] regs_23; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_23;
  reg [31:0] regs_24; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_24;
  reg [31:0] regs_25; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_25;
  reg [31:0] regs_26; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_26;
  reg [31:0] regs_27; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_27;
  reg [31:0] regs_28; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_28;
  reg [31:0] regs_29; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_29;
  reg [31:0] regs_30; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_30;
  reg [31:0] regs_31; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_31;
  reg [31:0] regs_32; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_32;
  reg [31:0] regs_33; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_33;
  reg [31:0] regs_34; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_34;
  reg [31:0] regs_35; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_35;
  reg [31:0] regs_36; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_36;
  reg [31:0] regs_37; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_37;
  reg [31:0] regs_38; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_38;
  reg [31:0] regs_39; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_39;
  reg [31:0] regs_40; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_40;
  reg [31:0] regs_41; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_41;
  reg [31:0] regs_42; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_42;
  reg [31:0] regs_43; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_43;
  reg [31:0] regs_44; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_44;
  reg [31:0] regs_45; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_45;
  reg [31:0] regs_46; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_46;
  reg [31:0] regs_47; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_47;
  reg [31:0] regs_48; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_48;
  reg [31:0] regs_49; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_49;
  reg [31:0] regs_50; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_50;
  reg [31:0] regs_51; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_51;
  reg [31:0] regs_52; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_52;
  reg [31:0] regs_53; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_53;
  reg [31:0] regs_54; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_54;
  reg [31:0] regs_55; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_55;
  reg [31:0] regs_56; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_56;
  reg [31:0] regs_57; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_57;
  reg [31:0] regs_58; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_58;
  reg [31:0] regs_59; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_59;
  reg [31:0] regs_60; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_60;
  reg [31:0] regs_61; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_61;
  reg [31:0] regs_62; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_62;
  reg [31:0] regs_63; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_63;
  reg [31:0] regs_64; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_64;
  reg [31:0] regs_65; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_65;
  reg [31:0] regs_66; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_66;
  reg [31:0] regs_67; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_67;
  reg [31:0] regs_68; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_68;
  reg [31:0] regs_69; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_69;
  reg [31:0] regs_70; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_70;
  reg [31:0] regs_71; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_71;
  reg [31:0] regs_72; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_72;
  reg [31:0] regs_73; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_73;
  reg [31:0] regs_74; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_74;
  reg [31:0] regs_75; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_75;
  reg [31:0] regs_76; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_76;
  reg [31:0] regs_77; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_77;
  reg [31:0] regs_78; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_78;
  reg [31:0] regs_79; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_79;
  reg [31:0] regs_80; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_80;
  reg [31:0] regs_81; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_81;
  reg [31:0] regs_82; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_82;
  reg [31:0] regs_83; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_83;
  reg [31:0] regs_84; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_84;
  reg [31:0] regs_85; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_85;
  reg [31:0] regs_86; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_86;
  reg [31:0] regs_87; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_87;
  reg [31:0] regs_88; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_88;
  reg [31:0] regs_89; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_89;
  reg [31:0] regs_90; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_90;
  reg [31:0] regs_91; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_91;
  reg [31:0] regs_92; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_92;
  reg [31:0] regs_93; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_93;
  reg [31:0] regs_94; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_94;
  reg [31:0] regs_95; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_95;
  reg [31:0] regs_96; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_96;
  reg [31:0] regs_97; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_97;
  reg [31:0] regs_98; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_98;
  reg [31:0] regs_99; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_99;
  reg [31:0] regs_100; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_100;
  reg [31:0] regs_101; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_101;
  reg [31:0] regs_102; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_102;
  reg [31:0] regs_103; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_103;
  reg [31:0] regs_104; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_104;
  reg [31:0] regs_105; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_105;
  reg [31:0] regs_106; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_106;
  reg [31:0] regs_107; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_107;
  reg [31:0] regs_108; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_108;
  reg [31:0] regs_109; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_109;
  reg [31:0] regs_110; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_110;
  reg [31:0] regs_111; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_111;
  reg [31:0] regs_112; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_112;
  reg [31:0] regs_113; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_113;
  reg [31:0] regs_114; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_114;
  reg [31:0] regs_115; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_115;
  reg [31:0] regs_116; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_116;
  reg [31:0] regs_117; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_117;
  reg [31:0] regs_118; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_118;
  reg [31:0] regs_119; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_119;
  reg [31:0] regs_120; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_120;
  reg [31:0] regs_121; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_121;
  reg [31:0] regs_122; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_122;
  reg [31:0] regs_123; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_123;
  reg [31:0] regs_124; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_124;
  reg [31:0] regs_125; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_125;
  reg [31:0] regs_126; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_126;
  reg [31:0] regs_127; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_127;
  reg [31:0] regs_128; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_128;
  reg [31:0] regs_129; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_129;
  reg [31:0] regs_130; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_130;
  reg [31:0] regs_131; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_131;
  reg [31:0] regs_132; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_132;
  reg [31:0] regs_133; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_133;
  reg [31:0] regs_134; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_134;
  reg [31:0] regs_135; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_135;
  reg [31:0] regs_136; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_136;
  reg [31:0] regs_137; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_137;
  reg [31:0] regs_138; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_138;
  reg [31:0] regs_139; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_139;
  reg [31:0] regs_140; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_140;
  reg [31:0] regs_141; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_141;
  reg [31:0] regs_142; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_142;
  reg [31:0] regs_143; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_143;
  reg [31:0] regs_144; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_144;
  reg [31:0] regs_145; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_145;
  reg [31:0] regs_146; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_146;
  reg [31:0] regs_147; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_147;
  reg [31:0] regs_148; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_148;
  reg [31:0] regs_149; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_149;
  reg [31:0] regs_150; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_150;
  reg [31:0] regs_151; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_151;
  reg [31:0] regs_152; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_152;
  reg [31:0] regs_153; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_153;
  reg [31:0] regs_154; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_154;
  reg [31:0] regs_155; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_155;
  reg [31:0] regs_156; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_156;
  reg [31:0] regs_157; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_157;
  reg [31:0] regs_158; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_158;
  reg [31:0] regs_159; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_159;
  reg [31:0] regs_160; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_160;
  reg [31:0] regs_161; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_161;
  reg [31:0] regs_162; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_162;
  reg [31:0] regs_163; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_163;
  reg [31:0] regs_164; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_164;
  reg [31:0] regs_165; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_165;
  reg [31:0] regs_166; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_166;
  reg [31:0] regs_167; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_167;
  reg [31:0] regs_168; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_168;
  reg [31:0] regs_169; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_169;
  reg [31:0] regs_170; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_170;
  reg [31:0] regs_171; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_171;
  reg [31:0] regs_172; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_172;
  reg [31:0] regs_173; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_173;
  reg [31:0] regs_174; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_174;
  reg [31:0] regs_175; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_175;
  reg [31:0] regs_176; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_176;
  reg [31:0] regs_177; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_177;
  reg [31:0] regs_178; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_178;
  reg [31:0] regs_179; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_179;
  reg [31:0] regs_180; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_180;
  reg [31:0] regs_181; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_181;
  reg [31:0] regs_182; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_182;
  reg [31:0] regs_183; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_183;
  reg [31:0] regs_184; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_184;
  reg [31:0] regs_185; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_185;
  reg [31:0] regs_186; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_186;
  reg [31:0] regs_187; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_187;
  reg [31:0] regs_188; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_188;
  reg [31:0] regs_189; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_189;
  reg [31:0] regs_190; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_190;
  reg [31:0] regs_191; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_191;
  reg [31:0] regs_192; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_192;
  reg [31:0] regs_193; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_193;
  reg [31:0] regs_194; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_194;
  reg [31:0] regs_195; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_195;
  reg [31:0] regs_196; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_196;
  reg [31:0] regs_197; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_197;
  reg [31:0] regs_198; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_198;
  reg [31:0] regs_199; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_199;
  reg [31:0] regs_200; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_200;
  reg [31:0] regs_201; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_201;
  reg [31:0] regs_202; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_202;
  reg [31:0] regs_203; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_203;
  reg [31:0] regs_204; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_204;
  reg [31:0] regs_205; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_205;
  reg [31:0] regs_206; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_206;
  reg [31:0] regs_207; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_207;
  reg [31:0] regs_208; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_208;
  reg [31:0] regs_209; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_209;
  assign io_out_bits_0_0 = regs_0; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_1 = regs_1; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_2 = regs_2; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_3 = regs_3; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_4 = regs_4; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_5 = regs_5; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_6 = regs_6; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_7 = regs_7; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_8 = regs_8; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_9 = regs_9; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_1_0 = regs_10; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_1_1 = regs_11; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_1_2 = regs_12; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_1_3 = regs_13; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_1_4 = regs_14; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_1_5 = regs_15; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_1_6 = regs_16; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_1_7 = regs_17; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_1_8 = regs_18; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_1_9 = regs_19; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_2_0 = regs_20; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_2_1 = regs_21; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_2_2 = regs_22; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_2_3 = regs_23; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_2_4 = regs_24; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_2_5 = regs_25; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_2_6 = regs_26; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_2_7 = regs_27; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_2_8 = regs_28; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_2_9 = regs_29; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_3_0 = regs_30; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_3_1 = regs_31; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_3_2 = regs_32; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_3_3 = regs_33; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_3_4 = regs_34; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_3_5 = regs_35; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_3_6 = regs_36; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_3_7 = regs_37; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_3_8 = regs_38; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_3_9 = regs_39; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_4_0 = regs_40; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_4_1 = regs_41; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_4_2 = regs_42; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_4_3 = regs_43; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_4_4 = regs_44; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_4_5 = regs_45; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_4_6 = regs_46; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_4_7 = regs_47; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_4_8 = regs_48; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_4_9 = regs_49; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_5_0 = regs_50; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_5_1 = regs_51; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_5_2 = regs_52; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_5_3 = regs_53; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_5_4 = regs_54; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_5_5 = regs_55; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_5_6 = regs_56; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_5_7 = regs_57; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_5_8 = regs_58; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_5_9 = regs_59; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_6_0 = regs_60; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_6_1 = regs_61; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_6_2 = regs_62; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_6_3 = regs_63; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_6_4 = regs_64; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_6_5 = regs_65; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_6_6 = regs_66; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_6_7 = regs_67; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_6_8 = regs_68; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_6_9 = regs_69; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_7_0 = regs_70; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_7_1 = regs_71; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_7_2 = regs_72; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_7_3 = regs_73; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_7_4 = regs_74; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_7_5 = regs_75; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_7_6 = regs_76; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_7_7 = regs_77; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_7_8 = regs_78; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_7_9 = regs_79; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_8_0 = regs_80; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_8_1 = regs_81; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_8_2 = regs_82; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_8_3 = regs_83; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_8_4 = regs_84; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_8_5 = regs_85; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_8_6 = regs_86; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_8_7 = regs_87; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_8_8 = regs_88; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_8_9 = regs_89; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_9_0 = regs_90; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_9_1 = regs_91; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_9_2 = regs_92; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_9_3 = regs_93; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_9_4 = regs_94; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_9_5 = regs_95; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_9_6 = regs_96; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_9_7 = regs_97; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_9_8 = regs_98; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_9_9 = regs_99; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_10_0 = regs_100; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_10_1 = regs_101; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_10_2 = regs_102; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_10_3 = regs_103; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_10_4 = regs_104; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_10_5 = regs_105; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_10_6 = regs_106; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_10_7 = regs_107; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_10_8 = regs_108; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_10_9 = regs_109; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_11_0 = regs_110; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_11_1 = regs_111; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_11_2 = regs_112; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_11_3 = regs_113; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_11_4 = regs_114; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_11_5 = regs_115; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_11_6 = regs_116; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_11_7 = regs_117; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_11_8 = regs_118; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_11_9 = regs_119; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_12_0 = regs_120; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_12_1 = regs_121; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_12_2 = regs_122; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_12_3 = regs_123; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_12_4 = regs_124; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_12_5 = regs_125; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_12_6 = regs_126; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_12_7 = regs_127; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_12_8 = regs_128; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_12_9 = regs_129; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_13_0 = regs_130; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_13_1 = regs_131; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_13_2 = regs_132; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_13_3 = regs_133; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_13_4 = regs_134; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_13_5 = regs_135; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_13_6 = regs_136; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_13_7 = regs_137; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_13_8 = regs_138; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_13_9 = regs_139; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_14_0 = regs_140; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_14_1 = regs_141; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_14_2 = regs_142; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_14_3 = regs_143; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_14_4 = regs_144; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_14_5 = regs_145; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_14_6 = regs_146; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_14_7 = regs_147; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_14_8 = regs_148; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_14_9 = regs_149; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_15_0 = regs_150; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_15_1 = regs_151; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_15_2 = regs_152; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_15_3 = regs_153; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_15_4 = regs_154; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_15_5 = regs_155; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_15_6 = regs_156; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_15_7 = regs_157; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_15_8 = regs_158; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_15_9 = regs_159; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_16_0 = regs_160; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_16_1 = regs_161; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_16_2 = regs_162; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_16_3 = regs_163; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_16_4 = regs_164; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_16_5 = regs_165; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_16_6 = regs_166; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_16_7 = regs_167; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_16_8 = regs_168; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_16_9 = regs_169; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_17_0 = regs_170; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_17_1 = regs_171; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_17_2 = regs_172; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_17_3 = regs_173; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_17_4 = regs_174; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_17_5 = regs_175; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_17_6 = regs_176; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_17_7 = regs_177; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_17_8 = regs_178; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_17_9 = regs_179; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_18_0 = regs_180; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_18_1 = regs_181; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_18_2 = regs_182; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_18_3 = regs_183; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_18_4 = regs_184; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_18_5 = regs_185; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_18_6 = regs_186; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_18_7 = regs_187; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_18_8 = regs_188; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_18_9 = regs_189; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_19_0 = regs_190; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_19_1 = regs_191; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_19_2 = regs_192; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_19_3 = regs_193; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_19_4 = regs_194; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_19_5 = regs_195; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_19_6 = regs_196; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_19_7 = regs_197; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_19_8 = regs_198; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_19_9 = regs_199; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_20_0 = regs_200; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_20_1 = regs_201; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_20_2 = regs_202; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_20_3 = regs_203; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_20_4 = regs_204; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_20_5 = regs_205; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_20_6 = regs_206; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_20_7 = regs_207; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_20_8 = regs_208; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_20_9 = regs_209; // @[MemoryBuffer.scala 65:25]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  regs_3 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  regs_4 = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  regs_5 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  regs_6 = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  regs_7 = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  regs_8 = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  regs_9 = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  regs_10 = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  regs_11 = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  regs_12 = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  regs_13 = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  regs_14 = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  regs_15 = _RAND_15[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  regs_16 = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  regs_17 = _RAND_17[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  regs_18 = _RAND_18[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  regs_19 = _RAND_19[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  regs_20 = _RAND_20[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  regs_21 = _RAND_21[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  regs_22 = _RAND_22[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  regs_23 = _RAND_23[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  regs_24 = _RAND_24[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  regs_25 = _RAND_25[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  regs_26 = _RAND_26[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  regs_27 = _RAND_27[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  regs_28 = _RAND_28[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  regs_29 = _RAND_29[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  regs_30 = _RAND_30[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  regs_31 = _RAND_31[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  regs_32 = _RAND_32[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  regs_33 = _RAND_33[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  regs_34 = _RAND_34[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  regs_35 = _RAND_35[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  regs_36 = _RAND_36[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  regs_37 = _RAND_37[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  regs_38 = _RAND_38[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  regs_39 = _RAND_39[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  regs_40 = _RAND_40[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  regs_41 = _RAND_41[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  regs_42 = _RAND_42[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  regs_43 = _RAND_43[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  regs_44 = _RAND_44[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  regs_45 = _RAND_45[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  regs_46 = _RAND_46[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  regs_47 = _RAND_47[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  regs_48 = _RAND_48[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  regs_49 = _RAND_49[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  regs_50 = _RAND_50[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  regs_51 = _RAND_51[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  regs_52 = _RAND_52[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  regs_53 = _RAND_53[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  regs_54 = _RAND_54[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  regs_55 = _RAND_55[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  regs_56 = _RAND_56[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  regs_57 = _RAND_57[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  regs_58 = _RAND_58[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  regs_59 = _RAND_59[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  regs_60 = _RAND_60[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  regs_61 = _RAND_61[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  regs_62 = _RAND_62[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  regs_63 = _RAND_63[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  regs_64 = _RAND_64[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  regs_65 = _RAND_65[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  regs_66 = _RAND_66[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  regs_67 = _RAND_67[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  regs_68 = _RAND_68[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  regs_69 = _RAND_69[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  regs_70 = _RAND_70[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  regs_71 = _RAND_71[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  regs_72 = _RAND_72[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  regs_73 = _RAND_73[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  regs_74 = _RAND_74[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  regs_75 = _RAND_75[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  regs_76 = _RAND_76[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  regs_77 = _RAND_77[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  regs_78 = _RAND_78[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  regs_79 = _RAND_79[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  regs_80 = _RAND_80[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  regs_81 = _RAND_81[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  regs_82 = _RAND_82[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  regs_83 = _RAND_83[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  regs_84 = _RAND_84[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  regs_85 = _RAND_85[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  regs_86 = _RAND_86[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  regs_87 = _RAND_87[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  regs_88 = _RAND_88[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  regs_89 = _RAND_89[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  regs_90 = _RAND_90[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  regs_91 = _RAND_91[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  regs_92 = _RAND_92[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  regs_93 = _RAND_93[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  regs_94 = _RAND_94[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  regs_95 = _RAND_95[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  regs_96 = _RAND_96[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  regs_97 = _RAND_97[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  regs_98 = _RAND_98[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  regs_99 = _RAND_99[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  regs_100 = _RAND_100[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  regs_101 = _RAND_101[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  regs_102 = _RAND_102[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  regs_103 = _RAND_103[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  regs_104 = _RAND_104[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  regs_105 = _RAND_105[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  regs_106 = _RAND_106[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  regs_107 = _RAND_107[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  regs_108 = _RAND_108[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  regs_109 = _RAND_109[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  regs_110 = _RAND_110[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  regs_111 = _RAND_111[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  regs_112 = _RAND_112[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  regs_113 = _RAND_113[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  regs_114 = _RAND_114[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  regs_115 = _RAND_115[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  regs_116 = _RAND_116[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  regs_117 = _RAND_117[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  regs_118 = _RAND_118[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  regs_119 = _RAND_119[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  regs_120 = _RAND_120[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  regs_121 = _RAND_121[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  regs_122 = _RAND_122[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  regs_123 = _RAND_123[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  regs_124 = _RAND_124[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  regs_125 = _RAND_125[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  regs_126 = _RAND_126[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  regs_127 = _RAND_127[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  regs_128 = _RAND_128[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  regs_129 = _RAND_129[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  regs_130 = _RAND_130[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  regs_131 = _RAND_131[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  regs_132 = _RAND_132[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  regs_133 = _RAND_133[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  regs_134 = _RAND_134[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  regs_135 = _RAND_135[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  regs_136 = _RAND_136[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  regs_137 = _RAND_137[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  regs_138 = _RAND_138[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  regs_139 = _RAND_139[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  regs_140 = _RAND_140[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  regs_141 = _RAND_141[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  regs_142 = _RAND_142[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  regs_143 = _RAND_143[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  regs_144 = _RAND_144[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  regs_145 = _RAND_145[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  regs_146 = _RAND_146[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{`RANDOM}};
  regs_147 = _RAND_147[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{`RANDOM}};
  regs_148 = _RAND_148[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{`RANDOM}};
  regs_149 = _RAND_149[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{`RANDOM}};
  regs_150 = _RAND_150[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{`RANDOM}};
  regs_151 = _RAND_151[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{`RANDOM}};
  regs_152 = _RAND_152[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  regs_153 = _RAND_153[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  regs_154 = _RAND_154[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  regs_155 = _RAND_155[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  regs_156 = _RAND_156[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  regs_157 = _RAND_157[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  regs_158 = _RAND_158[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  regs_159 = _RAND_159[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  regs_160 = _RAND_160[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  regs_161 = _RAND_161[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  regs_162 = _RAND_162[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  regs_163 = _RAND_163[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  regs_164 = _RAND_164[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  regs_165 = _RAND_165[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  regs_166 = _RAND_166[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  regs_167 = _RAND_167[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  regs_168 = _RAND_168[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{`RANDOM}};
  regs_169 = _RAND_169[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{`RANDOM}};
  regs_170 = _RAND_170[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  regs_171 = _RAND_171[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  regs_172 = _RAND_172[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{`RANDOM}};
  regs_173 = _RAND_173[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  regs_174 = _RAND_174[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  regs_175 = _RAND_175[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  regs_176 = _RAND_176[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  regs_177 = _RAND_177[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  regs_178 = _RAND_178[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{`RANDOM}};
  regs_179 = _RAND_179[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  regs_180 = _RAND_180[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{`RANDOM}};
  regs_181 = _RAND_181[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  regs_182 = _RAND_182[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  regs_183 = _RAND_183[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  regs_184 = _RAND_184[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  regs_185 = _RAND_185[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  regs_186 = _RAND_186[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  regs_187 = _RAND_187[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  regs_188 = _RAND_188[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{`RANDOM}};
  regs_189 = _RAND_189[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{`RANDOM}};
  regs_190 = _RAND_190[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{`RANDOM}};
  regs_191 = _RAND_191[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{`RANDOM}};
  regs_192 = _RAND_192[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{`RANDOM}};
  regs_193 = _RAND_193[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{`RANDOM}};
  regs_194 = _RAND_194[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{`RANDOM}};
  regs_195 = _RAND_195[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{`RANDOM}};
  regs_196 = _RAND_196[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{`RANDOM}};
  regs_197 = _RAND_197[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{`RANDOM}};
  regs_198 = _RAND_198[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{`RANDOM}};
  regs_199 = _RAND_199[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{`RANDOM}};
  regs_200 = _RAND_200[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{`RANDOM}};
  regs_201 = _RAND_201[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{`RANDOM}};
  regs_202 = _RAND_202[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{`RANDOM}};
  regs_203 = _RAND_203[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{`RANDOM}};
  regs_204 = _RAND_204[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{`RANDOM}};
  regs_205 = _RAND_205[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{`RANDOM}};
  regs_206 = _RAND_206[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{`RANDOM}};
  regs_207 = _RAND_207[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{`RANDOM}};
  regs_208 = _RAND_208[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{`RANDOM}};
  regs_209 = _RAND_209[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      regs_0 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_0 <= io_in_bits;
      end
    end
    if (reset) begin
      regs_1 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_1 <= regs_0;
      end
    end
    if (reset) begin
      regs_2 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_2 <= regs_1;
      end
    end
    if (reset) begin
      regs_3 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_3 <= regs_2;
      end
    end
    if (reset) begin
      regs_4 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_4 <= regs_3;
      end
    end
    if (reset) begin
      regs_5 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_5 <= regs_4;
      end
    end
    if (reset) begin
      regs_6 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_6 <= regs_5;
      end
    end
    if (reset) begin
      regs_7 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_7 <= regs_6;
      end
    end
    if (reset) begin
      regs_8 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_8 <= regs_7;
      end
    end
    if (reset) begin
      regs_9 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_9 <= regs_8;
      end
    end
    if (reset) begin
      regs_10 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_10 <= regs_9;
      end
    end
    if (reset) begin
      regs_11 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_11 <= regs_10;
      end
    end
    if (reset) begin
      regs_12 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_12 <= regs_11;
      end
    end
    if (reset) begin
      regs_13 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_13 <= regs_12;
      end
    end
    if (reset) begin
      regs_14 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_14 <= regs_13;
      end
    end
    if (reset) begin
      regs_15 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_15 <= regs_14;
      end
    end
    if (reset) begin
      regs_16 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_16 <= regs_15;
      end
    end
    if (reset) begin
      regs_17 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_17 <= regs_16;
      end
    end
    if (reset) begin
      regs_18 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_18 <= regs_17;
      end
    end
    if (reset) begin
      regs_19 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_19 <= regs_18;
      end
    end
    if (reset) begin
      regs_20 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_20 <= regs_19;
      end
    end
    if (reset) begin
      regs_21 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_21 <= regs_20;
      end
    end
    if (reset) begin
      regs_22 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_22 <= regs_21;
      end
    end
    if (reset) begin
      regs_23 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_23 <= regs_22;
      end
    end
    if (reset) begin
      regs_24 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_24 <= regs_23;
      end
    end
    if (reset) begin
      regs_25 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_25 <= regs_24;
      end
    end
    if (reset) begin
      regs_26 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_26 <= regs_25;
      end
    end
    if (reset) begin
      regs_27 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_27 <= regs_26;
      end
    end
    if (reset) begin
      regs_28 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_28 <= regs_27;
      end
    end
    if (reset) begin
      regs_29 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_29 <= regs_28;
      end
    end
    if (reset) begin
      regs_30 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_30 <= regs_29;
      end
    end
    if (reset) begin
      regs_31 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_31 <= regs_30;
      end
    end
    if (reset) begin
      regs_32 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_32 <= regs_31;
      end
    end
    if (reset) begin
      regs_33 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_33 <= regs_32;
      end
    end
    if (reset) begin
      regs_34 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_34 <= regs_33;
      end
    end
    if (reset) begin
      regs_35 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_35 <= regs_34;
      end
    end
    if (reset) begin
      regs_36 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_36 <= regs_35;
      end
    end
    if (reset) begin
      regs_37 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_37 <= regs_36;
      end
    end
    if (reset) begin
      regs_38 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_38 <= regs_37;
      end
    end
    if (reset) begin
      regs_39 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_39 <= regs_38;
      end
    end
    if (reset) begin
      regs_40 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_40 <= regs_39;
      end
    end
    if (reset) begin
      regs_41 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_41 <= regs_40;
      end
    end
    if (reset) begin
      regs_42 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_42 <= regs_41;
      end
    end
    if (reset) begin
      regs_43 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_43 <= regs_42;
      end
    end
    if (reset) begin
      regs_44 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_44 <= regs_43;
      end
    end
    if (reset) begin
      regs_45 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_45 <= regs_44;
      end
    end
    if (reset) begin
      regs_46 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_46 <= regs_45;
      end
    end
    if (reset) begin
      regs_47 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_47 <= regs_46;
      end
    end
    if (reset) begin
      regs_48 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_48 <= regs_47;
      end
    end
    if (reset) begin
      regs_49 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_49 <= regs_48;
      end
    end
    if (reset) begin
      regs_50 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_50 <= regs_49;
      end
    end
    if (reset) begin
      regs_51 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_51 <= regs_50;
      end
    end
    if (reset) begin
      regs_52 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_52 <= regs_51;
      end
    end
    if (reset) begin
      regs_53 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_53 <= regs_52;
      end
    end
    if (reset) begin
      regs_54 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_54 <= regs_53;
      end
    end
    if (reset) begin
      regs_55 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_55 <= regs_54;
      end
    end
    if (reset) begin
      regs_56 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_56 <= regs_55;
      end
    end
    if (reset) begin
      regs_57 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_57 <= regs_56;
      end
    end
    if (reset) begin
      regs_58 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_58 <= regs_57;
      end
    end
    if (reset) begin
      regs_59 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_59 <= regs_58;
      end
    end
    if (reset) begin
      regs_60 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_60 <= regs_59;
      end
    end
    if (reset) begin
      regs_61 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_61 <= regs_60;
      end
    end
    if (reset) begin
      regs_62 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_62 <= regs_61;
      end
    end
    if (reset) begin
      regs_63 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_63 <= regs_62;
      end
    end
    if (reset) begin
      regs_64 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_64 <= regs_63;
      end
    end
    if (reset) begin
      regs_65 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_65 <= regs_64;
      end
    end
    if (reset) begin
      regs_66 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_66 <= regs_65;
      end
    end
    if (reset) begin
      regs_67 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_67 <= regs_66;
      end
    end
    if (reset) begin
      regs_68 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_68 <= regs_67;
      end
    end
    if (reset) begin
      regs_69 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_69 <= regs_68;
      end
    end
    if (reset) begin
      regs_70 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_70 <= regs_69;
      end
    end
    if (reset) begin
      regs_71 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_71 <= regs_70;
      end
    end
    if (reset) begin
      regs_72 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_72 <= regs_71;
      end
    end
    if (reset) begin
      regs_73 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_73 <= regs_72;
      end
    end
    if (reset) begin
      regs_74 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_74 <= regs_73;
      end
    end
    if (reset) begin
      regs_75 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_75 <= regs_74;
      end
    end
    if (reset) begin
      regs_76 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_76 <= regs_75;
      end
    end
    if (reset) begin
      regs_77 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_77 <= regs_76;
      end
    end
    if (reset) begin
      regs_78 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_78 <= regs_77;
      end
    end
    if (reset) begin
      regs_79 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_79 <= regs_78;
      end
    end
    if (reset) begin
      regs_80 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_80 <= regs_79;
      end
    end
    if (reset) begin
      regs_81 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_81 <= regs_80;
      end
    end
    if (reset) begin
      regs_82 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_82 <= regs_81;
      end
    end
    if (reset) begin
      regs_83 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_83 <= regs_82;
      end
    end
    if (reset) begin
      regs_84 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_84 <= regs_83;
      end
    end
    if (reset) begin
      regs_85 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_85 <= regs_84;
      end
    end
    if (reset) begin
      regs_86 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_86 <= regs_85;
      end
    end
    if (reset) begin
      regs_87 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_87 <= regs_86;
      end
    end
    if (reset) begin
      regs_88 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_88 <= regs_87;
      end
    end
    if (reset) begin
      regs_89 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_89 <= regs_88;
      end
    end
    if (reset) begin
      regs_90 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_90 <= regs_89;
      end
    end
    if (reset) begin
      regs_91 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_91 <= regs_90;
      end
    end
    if (reset) begin
      regs_92 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_92 <= regs_91;
      end
    end
    if (reset) begin
      regs_93 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_93 <= regs_92;
      end
    end
    if (reset) begin
      regs_94 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_94 <= regs_93;
      end
    end
    if (reset) begin
      regs_95 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_95 <= regs_94;
      end
    end
    if (reset) begin
      regs_96 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_96 <= regs_95;
      end
    end
    if (reset) begin
      regs_97 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_97 <= regs_96;
      end
    end
    if (reset) begin
      regs_98 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_98 <= regs_97;
      end
    end
    if (reset) begin
      regs_99 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_99 <= regs_98;
      end
    end
    if (reset) begin
      regs_100 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_100 <= regs_99;
      end
    end
    if (reset) begin
      regs_101 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_101 <= regs_100;
      end
    end
    if (reset) begin
      regs_102 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_102 <= regs_101;
      end
    end
    if (reset) begin
      regs_103 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_103 <= regs_102;
      end
    end
    if (reset) begin
      regs_104 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_104 <= regs_103;
      end
    end
    if (reset) begin
      regs_105 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_105 <= regs_104;
      end
    end
    if (reset) begin
      regs_106 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_106 <= regs_105;
      end
    end
    if (reset) begin
      regs_107 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_107 <= regs_106;
      end
    end
    if (reset) begin
      regs_108 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_108 <= regs_107;
      end
    end
    if (reset) begin
      regs_109 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_109 <= regs_108;
      end
    end
    if (reset) begin
      regs_110 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_110 <= regs_109;
      end
    end
    if (reset) begin
      regs_111 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_111 <= regs_110;
      end
    end
    if (reset) begin
      regs_112 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_112 <= regs_111;
      end
    end
    if (reset) begin
      regs_113 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_113 <= regs_112;
      end
    end
    if (reset) begin
      regs_114 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_114 <= regs_113;
      end
    end
    if (reset) begin
      regs_115 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_115 <= regs_114;
      end
    end
    if (reset) begin
      regs_116 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_116 <= regs_115;
      end
    end
    if (reset) begin
      regs_117 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_117 <= regs_116;
      end
    end
    if (reset) begin
      regs_118 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_118 <= regs_117;
      end
    end
    if (reset) begin
      regs_119 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_119 <= regs_118;
      end
    end
    if (reset) begin
      regs_120 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_120 <= regs_119;
      end
    end
    if (reset) begin
      regs_121 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_121 <= regs_120;
      end
    end
    if (reset) begin
      regs_122 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_122 <= regs_121;
      end
    end
    if (reset) begin
      regs_123 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_123 <= regs_122;
      end
    end
    if (reset) begin
      regs_124 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_124 <= regs_123;
      end
    end
    if (reset) begin
      regs_125 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_125 <= regs_124;
      end
    end
    if (reset) begin
      regs_126 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_126 <= regs_125;
      end
    end
    if (reset) begin
      regs_127 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_127 <= regs_126;
      end
    end
    if (reset) begin
      regs_128 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_128 <= regs_127;
      end
    end
    if (reset) begin
      regs_129 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_129 <= regs_128;
      end
    end
    if (reset) begin
      regs_130 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_130 <= regs_129;
      end
    end
    if (reset) begin
      regs_131 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_131 <= regs_130;
      end
    end
    if (reset) begin
      regs_132 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_132 <= regs_131;
      end
    end
    if (reset) begin
      regs_133 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_133 <= regs_132;
      end
    end
    if (reset) begin
      regs_134 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_134 <= regs_133;
      end
    end
    if (reset) begin
      regs_135 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_135 <= regs_134;
      end
    end
    if (reset) begin
      regs_136 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_136 <= regs_135;
      end
    end
    if (reset) begin
      regs_137 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_137 <= regs_136;
      end
    end
    if (reset) begin
      regs_138 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_138 <= regs_137;
      end
    end
    if (reset) begin
      regs_139 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_139 <= regs_138;
      end
    end
    if (reset) begin
      regs_140 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_140 <= regs_139;
      end
    end
    if (reset) begin
      regs_141 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_141 <= regs_140;
      end
    end
    if (reset) begin
      regs_142 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_142 <= regs_141;
      end
    end
    if (reset) begin
      regs_143 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_143 <= regs_142;
      end
    end
    if (reset) begin
      regs_144 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_144 <= regs_143;
      end
    end
    if (reset) begin
      regs_145 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_145 <= regs_144;
      end
    end
    if (reset) begin
      regs_146 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_146 <= regs_145;
      end
    end
    if (reset) begin
      regs_147 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_147 <= regs_146;
      end
    end
    if (reset) begin
      regs_148 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_148 <= regs_147;
      end
    end
    if (reset) begin
      regs_149 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_149 <= regs_148;
      end
    end
    if (reset) begin
      regs_150 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_150 <= regs_149;
      end
    end
    if (reset) begin
      regs_151 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_151 <= regs_150;
      end
    end
    if (reset) begin
      regs_152 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_152 <= regs_151;
      end
    end
    if (reset) begin
      regs_153 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_153 <= regs_152;
      end
    end
    if (reset) begin
      regs_154 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_154 <= regs_153;
      end
    end
    if (reset) begin
      regs_155 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_155 <= regs_154;
      end
    end
    if (reset) begin
      regs_156 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_156 <= regs_155;
      end
    end
    if (reset) begin
      regs_157 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_157 <= regs_156;
      end
    end
    if (reset) begin
      regs_158 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_158 <= regs_157;
      end
    end
    if (reset) begin
      regs_159 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_159 <= regs_158;
      end
    end
    if (reset) begin
      regs_160 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_160 <= regs_159;
      end
    end
    if (reset) begin
      regs_161 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_161 <= regs_160;
      end
    end
    if (reset) begin
      regs_162 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_162 <= regs_161;
      end
    end
    if (reset) begin
      regs_163 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_163 <= regs_162;
      end
    end
    if (reset) begin
      regs_164 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_164 <= regs_163;
      end
    end
    if (reset) begin
      regs_165 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_165 <= regs_164;
      end
    end
    if (reset) begin
      regs_166 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_166 <= regs_165;
      end
    end
    if (reset) begin
      regs_167 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_167 <= regs_166;
      end
    end
    if (reset) begin
      regs_168 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_168 <= regs_167;
      end
    end
    if (reset) begin
      regs_169 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_169 <= regs_168;
      end
    end
    if (reset) begin
      regs_170 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_170 <= regs_169;
      end
    end
    if (reset) begin
      regs_171 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_171 <= regs_170;
      end
    end
    if (reset) begin
      regs_172 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_172 <= regs_171;
      end
    end
    if (reset) begin
      regs_173 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_173 <= regs_172;
      end
    end
    if (reset) begin
      regs_174 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_174 <= regs_173;
      end
    end
    if (reset) begin
      regs_175 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_175 <= regs_174;
      end
    end
    if (reset) begin
      regs_176 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_176 <= regs_175;
      end
    end
    if (reset) begin
      regs_177 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_177 <= regs_176;
      end
    end
    if (reset) begin
      regs_178 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_178 <= regs_177;
      end
    end
    if (reset) begin
      regs_179 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_179 <= regs_178;
      end
    end
    if (reset) begin
      regs_180 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_180 <= regs_179;
      end
    end
    if (reset) begin
      regs_181 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_181 <= regs_180;
      end
    end
    if (reset) begin
      regs_182 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_182 <= regs_181;
      end
    end
    if (reset) begin
      regs_183 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_183 <= regs_182;
      end
    end
    if (reset) begin
      regs_184 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_184 <= regs_183;
      end
    end
    if (reset) begin
      regs_185 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_185 <= regs_184;
      end
    end
    if (reset) begin
      regs_186 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_186 <= regs_185;
      end
    end
    if (reset) begin
      regs_187 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_187 <= regs_186;
      end
    end
    if (reset) begin
      regs_188 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_188 <= regs_187;
      end
    end
    if (reset) begin
      regs_189 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_189 <= regs_188;
      end
    end
    if (reset) begin
      regs_190 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_190 <= regs_189;
      end
    end
    if (reset) begin
      regs_191 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_191 <= regs_190;
      end
    end
    if (reset) begin
      regs_192 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_192 <= regs_191;
      end
    end
    if (reset) begin
      regs_193 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_193 <= regs_192;
      end
    end
    if (reset) begin
      regs_194 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_194 <= regs_193;
      end
    end
    if (reset) begin
      regs_195 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_195 <= regs_194;
      end
    end
    if (reset) begin
      regs_196 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_196 <= regs_195;
      end
    end
    if (reset) begin
      regs_197 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_197 <= regs_196;
      end
    end
    if (reset) begin
      regs_198 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_198 <= regs_197;
      end
    end
    if (reset) begin
      regs_199 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_199 <= regs_198;
      end
    end
    if (reset) begin
      regs_200 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_200 <= regs_199;
      end
    end
    if (reset) begin
      regs_201 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_201 <= regs_200;
      end
    end
    if (reset) begin
      regs_202 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_202 <= regs_201;
      end
    end
    if (reset) begin
      regs_203 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_203 <= regs_202;
      end
    end
    if (reset) begin
      regs_204 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_204 <= regs_203;
      end
    end
    if (reset) begin
      regs_205 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_205 <= regs_204;
      end
    end
    if (reset) begin
      regs_206 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_206 <= regs_205;
      end
    end
    if (reset) begin
      regs_207 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_207 <= regs_206;
      end
    end
    if (reset) begin
      regs_208 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_208 <= regs_207;
      end
    end
    if (reset) begin
      regs_209 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_209 <= regs_208;
      end
    end
  end
endmodule
module MemoryBuffer_2(
  input         clock,
  input         reset,
  input         io_in_valid,
  input  [31:0] io_in_bits,
  output [31:0] io_out_bits_0_0,
  output [31:0] io_out_bits_0_1,
  output [31:0] io_out_bits_0_2,
  output [31:0] io_out_bits_0_3,
  output [31:0] io_out_bits_0_4,
  output [31:0] io_out_bits_0_5,
  output [31:0] io_out_bits_0_6,
  output [31:0] io_out_bits_0_7,
  output [31:0] io_out_bits_0_8,
  output [31:0] io_out_bits_0_9,
  output [31:0] io_out_bits_1_0,
  output [31:0] io_out_bits_1_1,
  output [31:0] io_out_bits_1_2,
  output [31:0] io_out_bits_1_3,
  output [31:0] io_out_bits_1_4,
  output [31:0] io_out_bits_1_5,
  output [31:0] io_out_bits_1_6,
  output [31:0] io_out_bits_1_7,
  output [31:0] io_out_bits_1_8,
  output [31:0] io_out_bits_1_9,
  output [31:0] io_out_bits_2_0,
  output [31:0] io_out_bits_2_1,
  output [31:0] io_out_bits_2_2,
  output [31:0] io_out_bits_2_3,
  output [31:0] io_out_bits_2_4,
  output [31:0] io_out_bits_2_5,
  output [31:0] io_out_bits_2_6,
  output [31:0] io_out_bits_2_7,
  output [31:0] io_out_bits_2_8,
  output [31:0] io_out_bits_2_9
);
  reg [31:0] regs_0; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_0;
  reg [31:0] regs_1; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_1;
  reg [31:0] regs_2; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_2;
  reg [31:0] regs_3; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_3;
  reg [31:0] regs_4; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_4;
  reg [31:0] regs_5; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_5;
  reg [31:0] regs_6; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_6;
  reg [31:0] regs_7; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_7;
  reg [31:0] regs_8; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_8;
  reg [31:0] regs_9; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_9;
  reg [31:0] regs_10; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_10;
  reg [31:0] regs_11; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_11;
  reg [31:0] regs_12; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_12;
  reg [31:0] regs_13; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_13;
  reg [31:0] regs_14; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_14;
  reg [31:0] regs_15; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_15;
  reg [31:0] regs_16; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_16;
  reg [31:0] regs_17; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_17;
  reg [31:0] regs_18; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_18;
  reg [31:0] regs_19; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_19;
  reg [31:0] regs_20; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_20;
  reg [31:0] regs_21; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_21;
  reg [31:0] regs_22; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_22;
  reg [31:0] regs_23; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_23;
  reg [31:0] regs_24; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_24;
  reg [31:0] regs_25; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_25;
  reg [31:0] regs_26; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_26;
  reg [31:0] regs_27; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_27;
  reg [31:0] regs_28; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_28;
  reg [31:0] regs_29; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_29;
  assign io_out_bits_0_0 = regs_0; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_1 = regs_1; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_2 = regs_2; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_3 = regs_3; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_4 = regs_4; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_5 = regs_5; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_6 = regs_6; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_7 = regs_7; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_8 = regs_8; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_0_9 = regs_9; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_1_0 = regs_10; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_1_1 = regs_11; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_1_2 = regs_12; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_1_3 = regs_13; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_1_4 = regs_14; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_1_5 = regs_15; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_1_6 = regs_16; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_1_7 = regs_17; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_1_8 = regs_18; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_1_9 = regs_19; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_2_0 = regs_20; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_2_1 = regs_21; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_2_2 = regs_22; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_2_3 = regs_23; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_2_4 = regs_24; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_2_5 = regs_25; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_2_6 = regs_26; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_2_7 = regs_27; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_2_8 = regs_28; // @[MemoryBuffer.scala 65:25]
  assign io_out_bits_2_9 = regs_29; // @[MemoryBuffer.scala 65:25]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  regs_3 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  regs_4 = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  regs_5 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  regs_6 = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  regs_7 = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  regs_8 = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  regs_9 = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  regs_10 = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  regs_11 = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  regs_12 = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  regs_13 = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  regs_14 = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  regs_15 = _RAND_15[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  regs_16 = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  regs_17 = _RAND_17[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  regs_18 = _RAND_18[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  regs_19 = _RAND_19[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  regs_20 = _RAND_20[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  regs_21 = _RAND_21[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  regs_22 = _RAND_22[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  regs_23 = _RAND_23[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  regs_24 = _RAND_24[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  regs_25 = _RAND_25[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  regs_26 = _RAND_26[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  regs_27 = _RAND_27[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  regs_28 = _RAND_28[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  regs_29 = _RAND_29[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      regs_0 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_0 <= io_in_bits;
      end
    end
    if (reset) begin
      regs_1 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_1 <= regs_0;
      end
    end
    if (reset) begin
      regs_2 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_2 <= regs_1;
      end
    end
    if (reset) begin
      regs_3 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_3 <= regs_2;
      end
    end
    if (reset) begin
      regs_4 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_4 <= regs_3;
      end
    end
    if (reset) begin
      regs_5 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_5 <= regs_4;
      end
    end
    if (reset) begin
      regs_6 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_6 <= regs_5;
      end
    end
    if (reset) begin
      regs_7 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_7 <= regs_6;
      end
    end
    if (reset) begin
      regs_8 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_8 <= regs_7;
      end
    end
    if (reset) begin
      regs_9 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_9 <= regs_8;
      end
    end
    if (reset) begin
      regs_10 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_10 <= regs_9;
      end
    end
    if (reset) begin
      regs_11 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_11 <= regs_10;
      end
    end
    if (reset) begin
      regs_12 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_12 <= regs_11;
      end
    end
    if (reset) begin
      regs_13 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_13 <= regs_12;
      end
    end
    if (reset) begin
      regs_14 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_14 <= regs_13;
      end
    end
    if (reset) begin
      regs_15 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_15 <= regs_14;
      end
    end
    if (reset) begin
      regs_16 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_16 <= regs_15;
      end
    end
    if (reset) begin
      regs_17 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_17 <= regs_16;
      end
    end
    if (reset) begin
      regs_18 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_18 <= regs_17;
      end
    end
    if (reset) begin
      regs_19 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_19 <= regs_18;
      end
    end
    if (reset) begin
      regs_20 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_20 <= regs_19;
      end
    end
    if (reset) begin
      regs_21 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_21 <= regs_20;
      end
    end
    if (reset) begin
      regs_22 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_22 <= regs_21;
      end
    end
    if (reset) begin
      regs_23 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_23 <= regs_22;
      end
    end
    if (reset) begin
      regs_24 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_24 <= regs_23;
      end
    end
    if (reset) begin
      regs_25 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_25 <= regs_24;
      end
    end
    if (reset) begin
      regs_26 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_26 <= regs_25;
      end
    end
    if (reset) begin
      regs_27 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_27 <= regs_26;
      end
    end
    if (reset) begin
      regs_28 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_28 <= regs_27;
      end
    end
    if (reset) begin
      regs_29 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_29 <= regs_28;
      end
    end
  end
endmodule
module MemoryBuffer_3(
  input         clock,
  input         reset,
  input         io_in_valid,
  input  [31:0] io_in_bits,
  output [31:0] io_out_bits_0_0
);
  reg [31:0] regs_0; // @[MemoryBuffer.scala 39:21]
  reg [31:0] _RAND_0;
  assign io_out_bits_0_0 = regs_0; // @[MemoryBuffer.scala 65:25]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      regs_0 <= 32'sh0;
    end else begin
      if (io_in_valid) begin
        regs_0 <= io_in_bits;
      end
    end
  end
endmodule
module ConfigurationMemory(
  input         clock,
  input         reset,
  input         io_in_valid,
  input  [31:0] io_in_bits_wrdata,
  input  [2:0]  io_in_bits_wraddr,
  output [31:0] io_out_bits_confneuralNetsinputWeights_0_0,
  output [31:0] io_out_bits_confneuralNetsinputWeights_0_1,
  output [31:0] io_out_bits_confneuralNetsinputWeights_0_2,
  output [31:0] io_out_bits_confneuralNetsinputWeights_0_3,
  output [31:0] io_out_bits_confneuralNetsinputWeights_1_0,
  output [31:0] io_out_bits_confneuralNetsinputWeights_1_1,
  output [31:0] io_out_bits_confneuralNetsinputWeights_1_2,
  output [31:0] io_out_bits_confneuralNetsinputWeights_1_3,
  output [31:0] io_out_bits_confneuralNetsinputWeights_2_0,
  output [31:0] io_out_bits_confneuralNetsinputWeights_2_1,
  output [31:0] io_out_bits_confneuralNetsinputWeights_2_2,
  output [31:0] io_out_bits_confneuralNetsinputWeights_2_3,
  output [31:0] io_out_bits_confneuralNetsinputWeights_3_0,
  output [31:0] io_out_bits_confneuralNetsinputWeights_3_1,
  output [31:0] io_out_bits_confneuralNetsinputWeights_3_2,
  output [31:0] io_out_bits_confneuralNetsinputWeights_3_3,
  output [31:0] io_out_bits_confneuralNetsinputWeights_4_0,
  output [31:0] io_out_bits_confneuralNetsinputWeights_4_1,
  output [31:0] io_out_bits_confneuralNetsinputWeights_4_2,
  output [31:0] io_out_bits_confneuralNetsinputWeights_4_3,
  output [31:0] io_out_bits_confneuralNetsinputWeights_5_0,
  output [31:0] io_out_bits_confneuralNetsinputWeights_5_1,
  output [31:0] io_out_bits_confneuralNetsinputWeights_5_2,
  output [31:0] io_out_bits_confneuralNetsinputWeights_5_3,
  output [31:0] io_out_bits_confneuralNetsinputWeights_6_0,
  output [31:0] io_out_bits_confneuralNetsinputWeights_6_1,
  output [31:0] io_out_bits_confneuralNetsinputWeights_6_2,
  output [31:0] io_out_bits_confneuralNetsinputWeights_6_3,
  output [31:0] io_out_bits_confneuralNetsinputWeights_7_0,
  output [31:0] io_out_bits_confneuralNetsinputWeights_7_1,
  output [31:0] io_out_bits_confneuralNetsinputWeights_7_2,
  output [31:0] io_out_bits_confneuralNetsinputWeights_7_3,
  output [31:0] io_out_bits_confneuralNetsinputWeights_8_0,
  output [31:0] io_out_bits_confneuralNetsinputWeights_8_1,
  output [31:0] io_out_bits_confneuralNetsinputWeights_8_2,
  output [31:0] io_out_bits_confneuralNetsinputWeights_8_3,
  output [31:0] io_out_bits_confneuralNetsinputWeights_9_0,
  output [31:0] io_out_bits_confneuralNetsinputWeights_9_1,
  output [31:0] io_out_bits_confneuralNetsinputWeights_9_2,
  output [31:0] io_out_bits_confneuralNetsinputWeights_9_3,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_0_0,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_0_1,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_0_2,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_0_3,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_0_4,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_0_5,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_0_6,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_0_7,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_0_8,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_0_9,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_1_0,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_1_1,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_1_2,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_1_3,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_1_4,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_1_5,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_1_6,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_1_7,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_1_8,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_1_9,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_2_0,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_2_1,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_2_2,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_2_3,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_2_4,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_2_5,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_2_6,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_2_7,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_2_8,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_2_9,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_3_0,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_3_1,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_3_2,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_3_3,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_3_4,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_3_5,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_3_6,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_3_7,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_3_8,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_3_9,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_4_0,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_4_1,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_4_2,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_4_3,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_4_4,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_4_5,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_4_6,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_4_7,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_4_8,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_4_9,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_5_0,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_5_1,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_5_2,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_5_3,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_5_4,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_5_5,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_5_6,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_5_7,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_5_8,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_5_9,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_6_0,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_6_1,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_6_2,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_6_3,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_6_4,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_6_5,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_6_6,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_6_7,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_6_8,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_6_9,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_7_0,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_7_1,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_7_2,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_7_3,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_7_4,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_7_5,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_7_6,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_7_7,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_7_8,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_7_9,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_8_0,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_8_1,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_8_2,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_8_3,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_8_4,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_8_5,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_8_6,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_8_7,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_8_8,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_8_9,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_9_0,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_9_1,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_9_2,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_9_3,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_9_4,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_9_5,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_9_6,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_9_7,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_9_8,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_9_9,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_10_0,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_10_1,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_10_2,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_10_3,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_10_4,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_10_5,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_10_6,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_10_7,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_10_8,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_10_9,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_11_0,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_11_1,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_11_2,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_11_3,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_11_4,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_11_5,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_11_6,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_11_7,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_11_8,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_11_9,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_12_0,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_12_1,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_12_2,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_12_3,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_12_4,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_12_5,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_12_6,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_12_7,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_12_8,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_12_9,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_13_0,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_13_1,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_13_2,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_13_3,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_13_4,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_13_5,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_13_6,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_13_7,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_13_8,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_13_9,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_14_0,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_14_1,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_14_2,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_14_3,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_14_4,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_14_5,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_14_6,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_14_7,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_14_8,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_14_9,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_15_0,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_15_1,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_15_2,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_15_3,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_15_4,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_15_5,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_15_6,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_15_7,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_15_8,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_15_9,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_16_0,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_16_1,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_16_2,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_16_3,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_16_4,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_16_5,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_16_6,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_16_7,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_16_8,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_16_9,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_17_0,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_17_1,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_17_2,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_17_3,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_17_4,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_17_5,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_17_6,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_17_7,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_17_8,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_17_9,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_18_0,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_18_1,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_18_2,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_18_3,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_18_4,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_18_5,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_18_6,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_18_7,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_18_8,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_18_9,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_19_0,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_19_1,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_19_2,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_19_3,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_19_4,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_19_5,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_19_6,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_19_7,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_19_8,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_19_9,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_20_0,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_20_1,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_20_2,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_20_3,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_20_4,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_20_5,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_20_6,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_20_7,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_20_8,
  output [31:0] io_out_bits_confneuralNetsmidAndOutputWeights_20_9,
  output [31:0] io_out_bits_confneuralNetsbiasVecs_0_0,
  output [31:0] io_out_bits_confneuralNetsbiasVecs_0_1,
  output [31:0] io_out_bits_confneuralNetsbiasVecs_0_2,
  output [31:0] io_out_bits_confneuralNetsbiasVecs_0_3,
  output [31:0] io_out_bits_confneuralNetsbiasVecs_0_4,
  output [31:0] io_out_bits_confneuralNetsbiasVecs_0_5,
  output [31:0] io_out_bits_confneuralNetsbiasVecs_0_6,
  output [31:0] io_out_bits_confneuralNetsbiasVecs_0_7,
  output [31:0] io_out_bits_confneuralNetsbiasVecs_0_8,
  output [31:0] io_out_bits_confneuralNetsbiasVecs_0_9,
  output [31:0] io_out_bits_confneuralNetsbiasVecs_1_0,
  output [31:0] io_out_bits_confneuralNetsbiasVecs_1_1,
  output [31:0] io_out_bits_confneuralNetsbiasVecs_1_2,
  output [31:0] io_out_bits_confneuralNetsbiasVecs_1_3,
  output [31:0] io_out_bits_confneuralNetsbiasVecs_1_4,
  output [31:0] io_out_bits_confneuralNetsbiasVecs_1_5,
  output [31:0] io_out_bits_confneuralNetsbiasVecs_1_6,
  output [31:0] io_out_bits_confneuralNetsbiasVecs_1_7,
  output [31:0] io_out_bits_confneuralNetsbiasVecs_1_8,
  output [31:0] io_out_bits_confneuralNetsbiasVecs_1_9,
  output [31:0] io_out_bits_confneuralNetsbiasVecs_2_0,
  output [31:0] io_out_bits_confneuralNetsbiasVecs_2_1,
  output [31:0] io_out_bits_confneuralNetsbiasVecs_2_2,
  output [31:0] io_out_bits_confneuralNetsbiasVecs_2_3,
  output [31:0] io_out_bits_confneuralNetsbiasVecs_2_4,
  output [31:0] io_out_bits_confneuralNetsbiasVecs_2_5,
  output [31:0] io_out_bits_confneuralNetsbiasVecs_2_6,
  output [31:0] io_out_bits_confneuralNetsbiasVecs_2_7,
  output [31:0] io_out_bits_confneuralNetsbiasVecs_2_8,
  output [31:0] io_out_bits_confneuralNetsbiasVecs_2_9,
  output [31:0] io_out_bits_confneuralNetsoutputBias_0,
  output        io_out_bits_confInputMuxSel
);
  wire  neuralNetsinputWeightsMemory_clock; // @[ConfigurationMemory.scala 61:44]
  wire  neuralNetsinputWeightsMemory_reset; // @[ConfigurationMemory.scala 61:44]
  wire  neuralNetsinputWeightsMemory_io_in_valid; // @[ConfigurationMemory.scala 61:44]
  wire [31:0] neuralNetsinputWeightsMemory_io_in_bits; // @[ConfigurationMemory.scala 61:44]
  wire [31:0] neuralNetsinputWeightsMemory_io_out_bits_0_0; // @[ConfigurationMemory.scala 61:44]
  wire [31:0] neuralNetsinputWeightsMemory_io_out_bits_0_1; // @[ConfigurationMemory.scala 61:44]
  wire [31:0] neuralNetsinputWeightsMemory_io_out_bits_0_2; // @[ConfigurationMemory.scala 61:44]
  wire [31:0] neuralNetsinputWeightsMemory_io_out_bits_0_3; // @[ConfigurationMemory.scala 61:44]
  wire [31:0] neuralNetsinputWeightsMemory_io_out_bits_1_0; // @[ConfigurationMemory.scala 61:44]
  wire [31:0] neuralNetsinputWeightsMemory_io_out_bits_1_1; // @[ConfigurationMemory.scala 61:44]
  wire [31:0] neuralNetsinputWeightsMemory_io_out_bits_1_2; // @[ConfigurationMemory.scala 61:44]
  wire [31:0] neuralNetsinputWeightsMemory_io_out_bits_1_3; // @[ConfigurationMemory.scala 61:44]
  wire [31:0] neuralNetsinputWeightsMemory_io_out_bits_2_0; // @[ConfigurationMemory.scala 61:44]
  wire [31:0] neuralNetsinputWeightsMemory_io_out_bits_2_1; // @[ConfigurationMemory.scala 61:44]
  wire [31:0] neuralNetsinputWeightsMemory_io_out_bits_2_2; // @[ConfigurationMemory.scala 61:44]
  wire [31:0] neuralNetsinputWeightsMemory_io_out_bits_2_3; // @[ConfigurationMemory.scala 61:44]
  wire [31:0] neuralNetsinputWeightsMemory_io_out_bits_3_0; // @[ConfigurationMemory.scala 61:44]
  wire [31:0] neuralNetsinputWeightsMemory_io_out_bits_3_1; // @[ConfigurationMemory.scala 61:44]
  wire [31:0] neuralNetsinputWeightsMemory_io_out_bits_3_2; // @[ConfigurationMemory.scala 61:44]
  wire [31:0] neuralNetsinputWeightsMemory_io_out_bits_3_3; // @[ConfigurationMemory.scala 61:44]
  wire [31:0] neuralNetsinputWeightsMemory_io_out_bits_4_0; // @[ConfigurationMemory.scala 61:44]
  wire [31:0] neuralNetsinputWeightsMemory_io_out_bits_4_1; // @[ConfigurationMemory.scala 61:44]
  wire [31:0] neuralNetsinputWeightsMemory_io_out_bits_4_2; // @[ConfigurationMemory.scala 61:44]
  wire [31:0] neuralNetsinputWeightsMemory_io_out_bits_4_3; // @[ConfigurationMemory.scala 61:44]
  wire [31:0] neuralNetsinputWeightsMemory_io_out_bits_5_0; // @[ConfigurationMemory.scala 61:44]
  wire [31:0] neuralNetsinputWeightsMemory_io_out_bits_5_1; // @[ConfigurationMemory.scala 61:44]
  wire [31:0] neuralNetsinputWeightsMemory_io_out_bits_5_2; // @[ConfigurationMemory.scala 61:44]
  wire [31:0] neuralNetsinputWeightsMemory_io_out_bits_5_3; // @[ConfigurationMemory.scala 61:44]
  wire [31:0] neuralNetsinputWeightsMemory_io_out_bits_6_0; // @[ConfigurationMemory.scala 61:44]
  wire [31:0] neuralNetsinputWeightsMemory_io_out_bits_6_1; // @[ConfigurationMemory.scala 61:44]
  wire [31:0] neuralNetsinputWeightsMemory_io_out_bits_6_2; // @[ConfigurationMemory.scala 61:44]
  wire [31:0] neuralNetsinputWeightsMemory_io_out_bits_6_3; // @[ConfigurationMemory.scala 61:44]
  wire [31:0] neuralNetsinputWeightsMemory_io_out_bits_7_0; // @[ConfigurationMemory.scala 61:44]
  wire [31:0] neuralNetsinputWeightsMemory_io_out_bits_7_1; // @[ConfigurationMemory.scala 61:44]
  wire [31:0] neuralNetsinputWeightsMemory_io_out_bits_7_2; // @[ConfigurationMemory.scala 61:44]
  wire [31:0] neuralNetsinputWeightsMemory_io_out_bits_7_3; // @[ConfigurationMemory.scala 61:44]
  wire [31:0] neuralNetsinputWeightsMemory_io_out_bits_8_0; // @[ConfigurationMemory.scala 61:44]
  wire [31:0] neuralNetsinputWeightsMemory_io_out_bits_8_1; // @[ConfigurationMemory.scala 61:44]
  wire [31:0] neuralNetsinputWeightsMemory_io_out_bits_8_2; // @[ConfigurationMemory.scala 61:44]
  wire [31:0] neuralNetsinputWeightsMemory_io_out_bits_8_3; // @[ConfigurationMemory.scala 61:44]
  wire [31:0] neuralNetsinputWeightsMemory_io_out_bits_9_0; // @[ConfigurationMemory.scala 61:44]
  wire [31:0] neuralNetsinputWeightsMemory_io_out_bits_9_1; // @[ConfigurationMemory.scala 61:44]
  wire [31:0] neuralNetsinputWeightsMemory_io_out_bits_9_2; // @[ConfigurationMemory.scala 61:44]
  wire [31:0] neuralNetsinputWeightsMemory_io_out_bits_9_3; // @[ConfigurationMemory.scala 61:44]
  wire  neuralNetsmidAndOutputWeightsMemory_clock; // @[ConfigurationMemory.scala 73:51]
  wire  neuralNetsmidAndOutputWeightsMemory_reset; // @[ConfigurationMemory.scala 73:51]
  wire  neuralNetsmidAndOutputWeightsMemory_io_in_valid; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_in_bits; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_0_0; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_0_1; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_0_2; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_0_3; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_0_4; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_0_5; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_0_6; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_0_7; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_0_8; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_0_9; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_1_0; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_1_1; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_1_2; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_1_3; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_1_4; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_1_5; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_1_6; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_1_7; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_1_8; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_1_9; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_2_0; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_2_1; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_2_2; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_2_3; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_2_4; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_2_5; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_2_6; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_2_7; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_2_8; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_2_9; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_3_0; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_3_1; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_3_2; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_3_3; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_3_4; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_3_5; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_3_6; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_3_7; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_3_8; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_3_9; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_4_0; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_4_1; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_4_2; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_4_3; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_4_4; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_4_5; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_4_6; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_4_7; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_4_8; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_4_9; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_5_0; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_5_1; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_5_2; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_5_3; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_5_4; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_5_5; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_5_6; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_5_7; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_5_8; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_5_9; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_6_0; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_6_1; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_6_2; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_6_3; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_6_4; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_6_5; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_6_6; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_6_7; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_6_8; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_6_9; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_7_0; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_7_1; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_7_2; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_7_3; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_7_4; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_7_5; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_7_6; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_7_7; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_7_8; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_7_9; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_8_0; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_8_1; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_8_2; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_8_3; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_8_4; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_8_5; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_8_6; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_8_7; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_8_8; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_8_9; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_9_0; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_9_1; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_9_2; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_9_3; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_9_4; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_9_5; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_9_6; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_9_7; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_9_8; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_9_9; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_10_0; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_10_1; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_10_2; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_10_3; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_10_4; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_10_5; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_10_6; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_10_7; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_10_8; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_10_9; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_11_0; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_11_1; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_11_2; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_11_3; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_11_4; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_11_5; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_11_6; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_11_7; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_11_8; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_11_9; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_12_0; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_12_1; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_12_2; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_12_3; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_12_4; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_12_5; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_12_6; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_12_7; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_12_8; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_12_9; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_13_0; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_13_1; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_13_2; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_13_3; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_13_4; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_13_5; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_13_6; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_13_7; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_13_8; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_13_9; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_14_0; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_14_1; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_14_2; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_14_3; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_14_4; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_14_5; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_14_6; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_14_7; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_14_8; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_14_9; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_15_0; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_15_1; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_15_2; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_15_3; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_15_4; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_15_5; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_15_6; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_15_7; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_15_8; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_15_9; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_16_0; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_16_1; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_16_2; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_16_3; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_16_4; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_16_5; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_16_6; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_16_7; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_16_8; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_16_9; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_17_0; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_17_1; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_17_2; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_17_3; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_17_4; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_17_5; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_17_6; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_17_7; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_17_8; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_17_9; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_18_0; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_18_1; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_18_2; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_18_3; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_18_4; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_18_5; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_18_6; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_18_7; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_18_8; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_18_9; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_19_0; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_19_1; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_19_2; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_19_3; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_19_4; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_19_5; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_19_6; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_19_7; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_19_8; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_19_9; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_20_0; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_20_1; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_20_2; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_20_3; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_20_4; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_20_5; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_20_6; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_20_7; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_20_8; // @[ConfigurationMemory.scala 73:51]
  wire [31:0] neuralNetsmidAndOutputWeightsMemory_io_out_bits_20_9; // @[ConfigurationMemory.scala 73:51]
  wire  neuralNetsbiasVecsMemory_clock; // @[ConfigurationMemory.scala 84:40]
  wire  neuralNetsbiasVecsMemory_reset; // @[ConfigurationMemory.scala 84:40]
  wire  neuralNetsbiasVecsMemory_io_in_valid; // @[ConfigurationMemory.scala 84:40]
  wire [31:0] neuralNetsbiasVecsMemory_io_in_bits; // @[ConfigurationMemory.scala 84:40]
  wire [31:0] neuralNetsbiasVecsMemory_io_out_bits_0_0; // @[ConfigurationMemory.scala 84:40]
  wire [31:0] neuralNetsbiasVecsMemory_io_out_bits_0_1; // @[ConfigurationMemory.scala 84:40]
  wire [31:0] neuralNetsbiasVecsMemory_io_out_bits_0_2; // @[ConfigurationMemory.scala 84:40]
  wire [31:0] neuralNetsbiasVecsMemory_io_out_bits_0_3; // @[ConfigurationMemory.scala 84:40]
  wire [31:0] neuralNetsbiasVecsMemory_io_out_bits_0_4; // @[ConfigurationMemory.scala 84:40]
  wire [31:0] neuralNetsbiasVecsMemory_io_out_bits_0_5; // @[ConfigurationMemory.scala 84:40]
  wire [31:0] neuralNetsbiasVecsMemory_io_out_bits_0_6; // @[ConfigurationMemory.scala 84:40]
  wire [31:0] neuralNetsbiasVecsMemory_io_out_bits_0_7; // @[ConfigurationMemory.scala 84:40]
  wire [31:0] neuralNetsbiasVecsMemory_io_out_bits_0_8; // @[ConfigurationMemory.scala 84:40]
  wire [31:0] neuralNetsbiasVecsMemory_io_out_bits_0_9; // @[ConfigurationMemory.scala 84:40]
  wire [31:0] neuralNetsbiasVecsMemory_io_out_bits_1_0; // @[ConfigurationMemory.scala 84:40]
  wire [31:0] neuralNetsbiasVecsMemory_io_out_bits_1_1; // @[ConfigurationMemory.scala 84:40]
  wire [31:0] neuralNetsbiasVecsMemory_io_out_bits_1_2; // @[ConfigurationMemory.scala 84:40]
  wire [31:0] neuralNetsbiasVecsMemory_io_out_bits_1_3; // @[ConfigurationMemory.scala 84:40]
  wire [31:0] neuralNetsbiasVecsMemory_io_out_bits_1_4; // @[ConfigurationMemory.scala 84:40]
  wire [31:0] neuralNetsbiasVecsMemory_io_out_bits_1_5; // @[ConfigurationMemory.scala 84:40]
  wire [31:0] neuralNetsbiasVecsMemory_io_out_bits_1_6; // @[ConfigurationMemory.scala 84:40]
  wire [31:0] neuralNetsbiasVecsMemory_io_out_bits_1_7; // @[ConfigurationMemory.scala 84:40]
  wire [31:0] neuralNetsbiasVecsMemory_io_out_bits_1_8; // @[ConfigurationMemory.scala 84:40]
  wire [31:0] neuralNetsbiasVecsMemory_io_out_bits_1_9; // @[ConfigurationMemory.scala 84:40]
  wire [31:0] neuralNetsbiasVecsMemory_io_out_bits_2_0; // @[ConfigurationMemory.scala 84:40]
  wire [31:0] neuralNetsbiasVecsMemory_io_out_bits_2_1; // @[ConfigurationMemory.scala 84:40]
  wire [31:0] neuralNetsbiasVecsMemory_io_out_bits_2_2; // @[ConfigurationMemory.scala 84:40]
  wire [31:0] neuralNetsbiasVecsMemory_io_out_bits_2_3; // @[ConfigurationMemory.scala 84:40]
  wire [31:0] neuralNetsbiasVecsMemory_io_out_bits_2_4; // @[ConfigurationMemory.scala 84:40]
  wire [31:0] neuralNetsbiasVecsMemory_io_out_bits_2_5; // @[ConfigurationMemory.scala 84:40]
  wire [31:0] neuralNetsbiasVecsMemory_io_out_bits_2_6; // @[ConfigurationMemory.scala 84:40]
  wire [31:0] neuralNetsbiasVecsMemory_io_out_bits_2_7; // @[ConfigurationMemory.scala 84:40]
  wire [31:0] neuralNetsbiasVecsMemory_io_out_bits_2_8; // @[ConfigurationMemory.scala 84:40]
  wire [31:0] neuralNetsbiasVecsMemory_io_out_bits_2_9; // @[ConfigurationMemory.scala 84:40]
  wire  neuralNetsoutputBiasMemory_clock; // @[ConfigurationMemory.scala 96:42]
  wire  neuralNetsoutputBiasMemory_reset; // @[ConfigurationMemory.scala 96:42]
  wire  neuralNetsoutputBiasMemory_io_in_valid; // @[ConfigurationMemory.scala 96:42]
  wire [31:0] neuralNetsoutputBiasMemory_io_in_bits; // @[ConfigurationMemory.scala 96:42]
  wire [31:0] neuralNetsoutputBiasMemory_io_out_bits_0_0; // @[ConfigurationMemory.scala 96:42]
  wire  _T; // @[ConfigurationMemory.scala 64:68]
  wire  _T_2; // @[ConfigurationMemory.scala 76:75]
  wire  _T_4; // @[ConfigurationMemory.scala 87:64]
  wire  _T_6; // @[ConfigurationMemory.scala 99:66]
  reg  inputMuxSel; // @[ConfigurationMemory.scala 104:28]
  reg [31:0] _RAND_0;
  wire  _T_8; // @[ConfigurationMemory.scala 105:29]
  wire  _T_9; // @[ConfigurationMemory.scala 105:20]
  wire [31:0] _T_10; // @[ConfigurationMemory.scala 105:90]
  wire  _T_11; // @[ConfigurationMemory.scala 105:92]
  MemoryBuffer neuralNetsinputWeightsMemory ( // @[ConfigurationMemory.scala 61:44]
    .clock(neuralNetsinputWeightsMemory_clock),
    .reset(neuralNetsinputWeightsMemory_reset),
    .io_in_valid(neuralNetsinputWeightsMemory_io_in_valid),
    .io_in_bits(neuralNetsinputWeightsMemory_io_in_bits),
    .io_out_bits_0_0(neuralNetsinputWeightsMemory_io_out_bits_0_0),
    .io_out_bits_0_1(neuralNetsinputWeightsMemory_io_out_bits_0_1),
    .io_out_bits_0_2(neuralNetsinputWeightsMemory_io_out_bits_0_2),
    .io_out_bits_0_3(neuralNetsinputWeightsMemory_io_out_bits_0_3),
    .io_out_bits_1_0(neuralNetsinputWeightsMemory_io_out_bits_1_0),
    .io_out_bits_1_1(neuralNetsinputWeightsMemory_io_out_bits_1_1),
    .io_out_bits_1_2(neuralNetsinputWeightsMemory_io_out_bits_1_2),
    .io_out_bits_1_3(neuralNetsinputWeightsMemory_io_out_bits_1_3),
    .io_out_bits_2_0(neuralNetsinputWeightsMemory_io_out_bits_2_0),
    .io_out_bits_2_1(neuralNetsinputWeightsMemory_io_out_bits_2_1),
    .io_out_bits_2_2(neuralNetsinputWeightsMemory_io_out_bits_2_2),
    .io_out_bits_2_3(neuralNetsinputWeightsMemory_io_out_bits_2_3),
    .io_out_bits_3_0(neuralNetsinputWeightsMemory_io_out_bits_3_0),
    .io_out_bits_3_1(neuralNetsinputWeightsMemory_io_out_bits_3_1),
    .io_out_bits_3_2(neuralNetsinputWeightsMemory_io_out_bits_3_2),
    .io_out_bits_3_3(neuralNetsinputWeightsMemory_io_out_bits_3_3),
    .io_out_bits_4_0(neuralNetsinputWeightsMemory_io_out_bits_4_0),
    .io_out_bits_4_1(neuralNetsinputWeightsMemory_io_out_bits_4_1),
    .io_out_bits_4_2(neuralNetsinputWeightsMemory_io_out_bits_4_2),
    .io_out_bits_4_3(neuralNetsinputWeightsMemory_io_out_bits_4_3),
    .io_out_bits_5_0(neuralNetsinputWeightsMemory_io_out_bits_5_0),
    .io_out_bits_5_1(neuralNetsinputWeightsMemory_io_out_bits_5_1),
    .io_out_bits_5_2(neuralNetsinputWeightsMemory_io_out_bits_5_2),
    .io_out_bits_5_3(neuralNetsinputWeightsMemory_io_out_bits_5_3),
    .io_out_bits_6_0(neuralNetsinputWeightsMemory_io_out_bits_6_0),
    .io_out_bits_6_1(neuralNetsinputWeightsMemory_io_out_bits_6_1),
    .io_out_bits_6_2(neuralNetsinputWeightsMemory_io_out_bits_6_2),
    .io_out_bits_6_3(neuralNetsinputWeightsMemory_io_out_bits_6_3),
    .io_out_bits_7_0(neuralNetsinputWeightsMemory_io_out_bits_7_0),
    .io_out_bits_7_1(neuralNetsinputWeightsMemory_io_out_bits_7_1),
    .io_out_bits_7_2(neuralNetsinputWeightsMemory_io_out_bits_7_2),
    .io_out_bits_7_3(neuralNetsinputWeightsMemory_io_out_bits_7_3),
    .io_out_bits_8_0(neuralNetsinputWeightsMemory_io_out_bits_8_0),
    .io_out_bits_8_1(neuralNetsinputWeightsMemory_io_out_bits_8_1),
    .io_out_bits_8_2(neuralNetsinputWeightsMemory_io_out_bits_8_2),
    .io_out_bits_8_3(neuralNetsinputWeightsMemory_io_out_bits_8_3),
    .io_out_bits_9_0(neuralNetsinputWeightsMemory_io_out_bits_9_0),
    .io_out_bits_9_1(neuralNetsinputWeightsMemory_io_out_bits_9_1),
    .io_out_bits_9_2(neuralNetsinputWeightsMemory_io_out_bits_9_2),
    .io_out_bits_9_3(neuralNetsinputWeightsMemory_io_out_bits_9_3)
  );
  MemoryBuffer_1 neuralNetsmidAndOutputWeightsMemory ( // @[ConfigurationMemory.scala 73:51]
    .clock(neuralNetsmidAndOutputWeightsMemory_clock),
    .reset(neuralNetsmidAndOutputWeightsMemory_reset),
    .io_in_valid(neuralNetsmidAndOutputWeightsMemory_io_in_valid),
    .io_in_bits(neuralNetsmidAndOutputWeightsMemory_io_in_bits),
    .io_out_bits_0_0(neuralNetsmidAndOutputWeightsMemory_io_out_bits_0_0),
    .io_out_bits_0_1(neuralNetsmidAndOutputWeightsMemory_io_out_bits_0_1),
    .io_out_bits_0_2(neuralNetsmidAndOutputWeightsMemory_io_out_bits_0_2),
    .io_out_bits_0_3(neuralNetsmidAndOutputWeightsMemory_io_out_bits_0_3),
    .io_out_bits_0_4(neuralNetsmidAndOutputWeightsMemory_io_out_bits_0_4),
    .io_out_bits_0_5(neuralNetsmidAndOutputWeightsMemory_io_out_bits_0_5),
    .io_out_bits_0_6(neuralNetsmidAndOutputWeightsMemory_io_out_bits_0_6),
    .io_out_bits_0_7(neuralNetsmidAndOutputWeightsMemory_io_out_bits_0_7),
    .io_out_bits_0_8(neuralNetsmidAndOutputWeightsMemory_io_out_bits_0_8),
    .io_out_bits_0_9(neuralNetsmidAndOutputWeightsMemory_io_out_bits_0_9),
    .io_out_bits_1_0(neuralNetsmidAndOutputWeightsMemory_io_out_bits_1_0),
    .io_out_bits_1_1(neuralNetsmidAndOutputWeightsMemory_io_out_bits_1_1),
    .io_out_bits_1_2(neuralNetsmidAndOutputWeightsMemory_io_out_bits_1_2),
    .io_out_bits_1_3(neuralNetsmidAndOutputWeightsMemory_io_out_bits_1_3),
    .io_out_bits_1_4(neuralNetsmidAndOutputWeightsMemory_io_out_bits_1_4),
    .io_out_bits_1_5(neuralNetsmidAndOutputWeightsMemory_io_out_bits_1_5),
    .io_out_bits_1_6(neuralNetsmidAndOutputWeightsMemory_io_out_bits_1_6),
    .io_out_bits_1_7(neuralNetsmidAndOutputWeightsMemory_io_out_bits_1_7),
    .io_out_bits_1_8(neuralNetsmidAndOutputWeightsMemory_io_out_bits_1_8),
    .io_out_bits_1_9(neuralNetsmidAndOutputWeightsMemory_io_out_bits_1_9),
    .io_out_bits_2_0(neuralNetsmidAndOutputWeightsMemory_io_out_bits_2_0),
    .io_out_bits_2_1(neuralNetsmidAndOutputWeightsMemory_io_out_bits_2_1),
    .io_out_bits_2_2(neuralNetsmidAndOutputWeightsMemory_io_out_bits_2_2),
    .io_out_bits_2_3(neuralNetsmidAndOutputWeightsMemory_io_out_bits_2_3),
    .io_out_bits_2_4(neuralNetsmidAndOutputWeightsMemory_io_out_bits_2_4),
    .io_out_bits_2_5(neuralNetsmidAndOutputWeightsMemory_io_out_bits_2_5),
    .io_out_bits_2_6(neuralNetsmidAndOutputWeightsMemory_io_out_bits_2_6),
    .io_out_bits_2_7(neuralNetsmidAndOutputWeightsMemory_io_out_bits_2_7),
    .io_out_bits_2_8(neuralNetsmidAndOutputWeightsMemory_io_out_bits_2_8),
    .io_out_bits_2_9(neuralNetsmidAndOutputWeightsMemory_io_out_bits_2_9),
    .io_out_bits_3_0(neuralNetsmidAndOutputWeightsMemory_io_out_bits_3_0),
    .io_out_bits_3_1(neuralNetsmidAndOutputWeightsMemory_io_out_bits_3_1),
    .io_out_bits_3_2(neuralNetsmidAndOutputWeightsMemory_io_out_bits_3_2),
    .io_out_bits_3_3(neuralNetsmidAndOutputWeightsMemory_io_out_bits_3_3),
    .io_out_bits_3_4(neuralNetsmidAndOutputWeightsMemory_io_out_bits_3_4),
    .io_out_bits_3_5(neuralNetsmidAndOutputWeightsMemory_io_out_bits_3_5),
    .io_out_bits_3_6(neuralNetsmidAndOutputWeightsMemory_io_out_bits_3_6),
    .io_out_bits_3_7(neuralNetsmidAndOutputWeightsMemory_io_out_bits_3_7),
    .io_out_bits_3_8(neuralNetsmidAndOutputWeightsMemory_io_out_bits_3_8),
    .io_out_bits_3_9(neuralNetsmidAndOutputWeightsMemory_io_out_bits_3_9),
    .io_out_bits_4_0(neuralNetsmidAndOutputWeightsMemory_io_out_bits_4_0),
    .io_out_bits_4_1(neuralNetsmidAndOutputWeightsMemory_io_out_bits_4_1),
    .io_out_bits_4_2(neuralNetsmidAndOutputWeightsMemory_io_out_bits_4_2),
    .io_out_bits_4_3(neuralNetsmidAndOutputWeightsMemory_io_out_bits_4_3),
    .io_out_bits_4_4(neuralNetsmidAndOutputWeightsMemory_io_out_bits_4_4),
    .io_out_bits_4_5(neuralNetsmidAndOutputWeightsMemory_io_out_bits_4_5),
    .io_out_bits_4_6(neuralNetsmidAndOutputWeightsMemory_io_out_bits_4_6),
    .io_out_bits_4_7(neuralNetsmidAndOutputWeightsMemory_io_out_bits_4_7),
    .io_out_bits_4_8(neuralNetsmidAndOutputWeightsMemory_io_out_bits_4_8),
    .io_out_bits_4_9(neuralNetsmidAndOutputWeightsMemory_io_out_bits_4_9),
    .io_out_bits_5_0(neuralNetsmidAndOutputWeightsMemory_io_out_bits_5_0),
    .io_out_bits_5_1(neuralNetsmidAndOutputWeightsMemory_io_out_bits_5_1),
    .io_out_bits_5_2(neuralNetsmidAndOutputWeightsMemory_io_out_bits_5_2),
    .io_out_bits_5_3(neuralNetsmidAndOutputWeightsMemory_io_out_bits_5_3),
    .io_out_bits_5_4(neuralNetsmidAndOutputWeightsMemory_io_out_bits_5_4),
    .io_out_bits_5_5(neuralNetsmidAndOutputWeightsMemory_io_out_bits_5_5),
    .io_out_bits_5_6(neuralNetsmidAndOutputWeightsMemory_io_out_bits_5_6),
    .io_out_bits_5_7(neuralNetsmidAndOutputWeightsMemory_io_out_bits_5_7),
    .io_out_bits_5_8(neuralNetsmidAndOutputWeightsMemory_io_out_bits_5_8),
    .io_out_bits_5_9(neuralNetsmidAndOutputWeightsMemory_io_out_bits_5_9),
    .io_out_bits_6_0(neuralNetsmidAndOutputWeightsMemory_io_out_bits_6_0),
    .io_out_bits_6_1(neuralNetsmidAndOutputWeightsMemory_io_out_bits_6_1),
    .io_out_bits_6_2(neuralNetsmidAndOutputWeightsMemory_io_out_bits_6_2),
    .io_out_bits_6_3(neuralNetsmidAndOutputWeightsMemory_io_out_bits_6_3),
    .io_out_bits_6_4(neuralNetsmidAndOutputWeightsMemory_io_out_bits_6_4),
    .io_out_bits_6_5(neuralNetsmidAndOutputWeightsMemory_io_out_bits_6_5),
    .io_out_bits_6_6(neuralNetsmidAndOutputWeightsMemory_io_out_bits_6_6),
    .io_out_bits_6_7(neuralNetsmidAndOutputWeightsMemory_io_out_bits_6_7),
    .io_out_bits_6_8(neuralNetsmidAndOutputWeightsMemory_io_out_bits_6_8),
    .io_out_bits_6_9(neuralNetsmidAndOutputWeightsMemory_io_out_bits_6_9),
    .io_out_bits_7_0(neuralNetsmidAndOutputWeightsMemory_io_out_bits_7_0),
    .io_out_bits_7_1(neuralNetsmidAndOutputWeightsMemory_io_out_bits_7_1),
    .io_out_bits_7_2(neuralNetsmidAndOutputWeightsMemory_io_out_bits_7_2),
    .io_out_bits_7_3(neuralNetsmidAndOutputWeightsMemory_io_out_bits_7_3),
    .io_out_bits_7_4(neuralNetsmidAndOutputWeightsMemory_io_out_bits_7_4),
    .io_out_bits_7_5(neuralNetsmidAndOutputWeightsMemory_io_out_bits_7_5),
    .io_out_bits_7_6(neuralNetsmidAndOutputWeightsMemory_io_out_bits_7_6),
    .io_out_bits_7_7(neuralNetsmidAndOutputWeightsMemory_io_out_bits_7_7),
    .io_out_bits_7_8(neuralNetsmidAndOutputWeightsMemory_io_out_bits_7_8),
    .io_out_bits_7_9(neuralNetsmidAndOutputWeightsMemory_io_out_bits_7_9),
    .io_out_bits_8_0(neuralNetsmidAndOutputWeightsMemory_io_out_bits_8_0),
    .io_out_bits_8_1(neuralNetsmidAndOutputWeightsMemory_io_out_bits_8_1),
    .io_out_bits_8_2(neuralNetsmidAndOutputWeightsMemory_io_out_bits_8_2),
    .io_out_bits_8_3(neuralNetsmidAndOutputWeightsMemory_io_out_bits_8_3),
    .io_out_bits_8_4(neuralNetsmidAndOutputWeightsMemory_io_out_bits_8_4),
    .io_out_bits_8_5(neuralNetsmidAndOutputWeightsMemory_io_out_bits_8_5),
    .io_out_bits_8_6(neuralNetsmidAndOutputWeightsMemory_io_out_bits_8_6),
    .io_out_bits_8_7(neuralNetsmidAndOutputWeightsMemory_io_out_bits_8_7),
    .io_out_bits_8_8(neuralNetsmidAndOutputWeightsMemory_io_out_bits_8_8),
    .io_out_bits_8_9(neuralNetsmidAndOutputWeightsMemory_io_out_bits_8_9),
    .io_out_bits_9_0(neuralNetsmidAndOutputWeightsMemory_io_out_bits_9_0),
    .io_out_bits_9_1(neuralNetsmidAndOutputWeightsMemory_io_out_bits_9_1),
    .io_out_bits_9_2(neuralNetsmidAndOutputWeightsMemory_io_out_bits_9_2),
    .io_out_bits_9_3(neuralNetsmidAndOutputWeightsMemory_io_out_bits_9_3),
    .io_out_bits_9_4(neuralNetsmidAndOutputWeightsMemory_io_out_bits_9_4),
    .io_out_bits_9_5(neuralNetsmidAndOutputWeightsMemory_io_out_bits_9_5),
    .io_out_bits_9_6(neuralNetsmidAndOutputWeightsMemory_io_out_bits_9_6),
    .io_out_bits_9_7(neuralNetsmidAndOutputWeightsMemory_io_out_bits_9_7),
    .io_out_bits_9_8(neuralNetsmidAndOutputWeightsMemory_io_out_bits_9_8),
    .io_out_bits_9_9(neuralNetsmidAndOutputWeightsMemory_io_out_bits_9_9),
    .io_out_bits_10_0(neuralNetsmidAndOutputWeightsMemory_io_out_bits_10_0),
    .io_out_bits_10_1(neuralNetsmidAndOutputWeightsMemory_io_out_bits_10_1),
    .io_out_bits_10_2(neuralNetsmidAndOutputWeightsMemory_io_out_bits_10_2),
    .io_out_bits_10_3(neuralNetsmidAndOutputWeightsMemory_io_out_bits_10_3),
    .io_out_bits_10_4(neuralNetsmidAndOutputWeightsMemory_io_out_bits_10_4),
    .io_out_bits_10_5(neuralNetsmidAndOutputWeightsMemory_io_out_bits_10_5),
    .io_out_bits_10_6(neuralNetsmidAndOutputWeightsMemory_io_out_bits_10_6),
    .io_out_bits_10_7(neuralNetsmidAndOutputWeightsMemory_io_out_bits_10_7),
    .io_out_bits_10_8(neuralNetsmidAndOutputWeightsMemory_io_out_bits_10_8),
    .io_out_bits_10_9(neuralNetsmidAndOutputWeightsMemory_io_out_bits_10_9),
    .io_out_bits_11_0(neuralNetsmidAndOutputWeightsMemory_io_out_bits_11_0),
    .io_out_bits_11_1(neuralNetsmidAndOutputWeightsMemory_io_out_bits_11_1),
    .io_out_bits_11_2(neuralNetsmidAndOutputWeightsMemory_io_out_bits_11_2),
    .io_out_bits_11_3(neuralNetsmidAndOutputWeightsMemory_io_out_bits_11_3),
    .io_out_bits_11_4(neuralNetsmidAndOutputWeightsMemory_io_out_bits_11_4),
    .io_out_bits_11_5(neuralNetsmidAndOutputWeightsMemory_io_out_bits_11_5),
    .io_out_bits_11_6(neuralNetsmidAndOutputWeightsMemory_io_out_bits_11_6),
    .io_out_bits_11_7(neuralNetsmidAndOutputWeightsMemory_io_out_bits_11_7),
    .io_out_bits_11_8(neuralNetsmidAndOutputWeightsMemory_io_out_bits_11_8),
    .io_out_bits_11_9(neuralNetsmidAndOutputWeightsMemory_io_out_bits_11_9),
    .io_out_bits_12_0(neuralNetsmidAndOutputWeightsMemory_io_out_bits_12_0),
    .io_out_bits_12_1(neuralNetsmidAndOutputWeightsMemory_io_out_bits_12_1),
    .io_out_bits_12_2(neuralNetsmidAndOutputWeightsMemory_io_out_bits_12_2),
    .io_out_bits_12_3(neuralNetsmidAndOutputWeightsMemory_io_out_bits_12_3),
    .io_out_bits_12_4(neuralNetsmidAndOutputWeightsMemory_io_out_bits_12_4),
    .io_out_bits_12_5(neuralNetsmidAndOutputWeightsMemory_io_out_bits_12_5),
    .io_out_bits_12_6(neuralNetsmidAndOutputWeightsMemory_io_out_bits_12_6),
    .io_out_bits_12_7(neuralNetsmidAndOutputWeightsMemory_io_out_bits_12_7),
    .io_out_bits_12_8(neuralNetsmidAndOutputWeightsMemory_io_out_bits_12_8),
    .io_out_bits_12_9(neuralNetsmidAndOutputWeightsMemory_io_out_bits_12_9),
    .io_out_bits_13_0(neuralNetsmidAndOutputWeightsMemory_io_out_bits_13_0),
    .io_out_bits_13_1(neuralNetsmidAndOutputWeightsMemory_io_out_bits_13_1),
    .io_out_bits_13_2(neuralNetsmidAndOutputWeightsMemory_io_out_bits_13_2),
    .io_out_bits_13_3(neuralNetsmidAndOutputWeightsMemory_io_out_bits_13_3),
    .io_out_bits_13_4(neuralNetsmidAndOutputWeightsMemory_io_out_bits_13_4),
    .io_out_bits_13_5(neuralNetsmidAndOutputWeightsMemory_io_out_bits_13_5),
    .io_out_bits_13_6(neuralNetsmidAndOutputWeightsMemory_io_out_bits_13_6),
    .io_out_bits_13_7(neuralNetsmidAndOutputWeightsMemory_io_out_bits_13_7),
    .io_out_bits_13_8(neuralNetsmidAndOutputWeightsMemory_io_out_bits_13_8),
    .io_out_bits_13_9(neuralNetsmidAndOutputWeightsMemory_io_out_bits_13_9),
    .io_out_bits_14_0(neuralNetsmidAndOutputWeightsMemory_io_out_bits_14_0),
    .io_out_bits_14_1(neuralNetsmidAndOutputWeightsMemory_io_out_bits_14_1),
    .io_out_bits_14_2(neuralNetsmidAndOutputWeightsMemory_io_out_bits_14_2),
    .io_out_bits_14_3(neuralNetsmidAndOutputWeightsMemory_io_out_bits_14_3),
    .io_out_bits_14_4(neuralNetsmidAndOutputWeightsMemory_io_out_bits_14_4),
    .io_out_bits_14_5(neuralNetsmidAndOutputWeightsMemory_io_out_bits_14_5),
    .io_out_bits_14_6(neuralNetsmidAndOutputWeightsMemory_io_out_bits_14_6),
    .io_out_bits_14_7(neuralNetsmidAndOutputWeightsMemory_io_out_bits_14_7),
    .io_out_bits_14_8(neuralNetsmidAndOutputWeightsMemory_io_out_bits_14_8),
    .io_out_bits_14_9(neuralNetsmidAndOutputWeightsMemory_io_out_bits_14_9),
    .io_out_bits_15_0(neuralNetsmidAndOutputWeightsMemory_io_out_bits_15_0),
    .io_out_bits_15_1(neuralNetsmidAndOutputWeightsMemory_io_out_bits_15_1),
    .io_out_bits_15_2(neuralNetsmidAndOutputWeightsMemory_io_out_bits_15_2),
    .io_out_bits_15_3(neuralNetsmidAndOutputWeightsMemory_io_out_bits_15_3),
    .io_out_bits_15_4(neuralNetsmidAndOutputWeightsMemory_io_out_bits_15_4),
    .io_out_bits_15_5(neuralNetsmidAndOutputWeightsMemory_io_out_bits_15_5),
    .io_out_bits_15_6(neuralNetsmidAndOutputWeightsMemory_io_out_bits_15_6),
    .io_out_bits_15_7(neuralNetsmidAndOutputWeightsMemory_io_out_bits_15_7),
    .io_out_bits_15_8(neuralNetsmidAndOutputWeightsMemory_io_out_bits_15_8),
    .io_out_bits_15_9(neuralNetsmidAndOutputWeightsMemory_io_out_bits_15_9),
    .io_out_bits_16_0(neuralNetsmidAndOutputWeightsMemory_io_out_bits_16_0),
    .io_out_bits_16_1(neuralNetsmidAndOutputWeightsMemory_io_out_bits_16_1),
    .io_out_bits_16_2(neuralNetsmidAndOutputWeightsMemory_io_out_bits_16_2),
    .io_out_bits_16_3(neuralNetsmidAndOutputWeightsMemory_io_out_bits_16_3),
    .io_out_bits_16_4(neuralNetsmidAndOutputWeightsMemory_io_out_bits_16_4),
    .io_out_bits_16_5(neuralNetsmidAndOutputWeightsMemory_io_out_bits_16_5),
    .io_out_bits_16_6(neuralNetsmidAndOutputWeightsMemory_io_out_bits_16_6),
    .io_out_bits_16_7(neuralNetsmidAndOutputWeightsMemory_io_out_bits_16_7),
    .io_out_bits_16_8(neuralNetsmidAndOutputWeightsMemory_io_out_bits_16_8),
    .io_out_bits_16_9(neuralNetsmidAndOutputWeightsMemory_io_out_bits_16_9),
    .io_out_bits_17_0(neuralNetsmidAndOutputWeightsMemory_io_out_bits_17_0),
    .io_out_bits_17_1(neuralNetsmidAndOutputWeightsMemory_io_out_bits_17_1),
    .io_out_bits_17_2(neuralNetsmidAndOutputWeightsMemory_io_out_bits_17_2),
    .io_out_bits_17_3(neuralNetsmidAndOutputWeightsMemory_io_out_bits_17_3),
    .io_out_bits_17_4(neuralNetsmidAndOutputWeightsMemory_io_out_bits_17_4),
    .io_out_bits_17_5(neuralNetsmidAndOutputWeightsMemory_io_out_bits_17_5),
    .io_out_bits_17_6(neuralNetsmidAndOutputWeightsMemory_io_out_bits_17_6),
    .io_out_bits_17_7(neuralNetsmidAndOutputWeightsMemory_io_out_bits_17_7),
    .io_out_bits_17_8(neuralNetsmidAndOutputWeightsMemory_io_out_bits_17_8),
    .io_out_bits_17_9(neuralNetsmidAndOutputWeightsMemory_io_out_bits_17_9),
    .io_out_bits_18_0(neuralNetsmidAndOutputWeightsMemory_io_out_bits_18_0),
    .io_out_bits_18_1(neuralNetsmidAndOutputWeightsMemory_io_out_bits_18_1),
    .io_out_bits_18_2(neuralNetsmidAndOutputWeightsMemory_io_out_bits_18_2),
    .io_out_bits_18_3(neuralNetsmidAndOutputWeightsMemory_io_out_bits_18_3),
    .io_out_bits_18_4(neuralNetsmidAndOutputWeightsMemory_io_out_bits_18_4),
    .io_out_bits_18_5(neuralNetsmidAndOutputWeightsMemory_io_out_bits_18_5),
    .io_out_bits_18_6(neuralNetsmidAndOutputWeightsMemory_io_out_bits_18_6),
    .io_out_bits_18_7(neuralNetsmidAndOutputWeightsMemory_io_out_bits_18_7),
    .io_out_bits_18_8(neuralNetsmidAndOutputWeightsMemory_io_out_bits_18_8),
    .io_out_bits_18_9(neuralNetsmidAndOutputWeightsMemory_io_out_bits_18_9),
    .io_out_bits_19_0(neuralNetsmidAndOutputWeightsMemory_io_out_bits_19_0),
    .io_out_bits_19_1(neuralNetsmidAndOutputWeightsMemory_io_out_bits_19_1),
    .io_out_bits_19_2(neuralNetsmidAndOutputWeightsMemory_io_out_bits_19_2),
    .io_out_bits_19_3(neuralNetsmidAndOutputWeightsMemory_io_out_bits_19_3),
    .io_out_bits_19_4(neuralNetsmidAndOutputWeightsMemory_io_out_bits_19_4),
    .io_out_bits_19_5(neuralNetsmidAndOutputWeightsMemory_io_out_bits_19_5),
    .io_out_bits_19_6(neuralNetsmidAndOutputWeightsMemory_io_out_bits_19_6),
    .io_out_bits_19_7(neuralNetsmidAndOutputWeightsMemory_io_out_bits_19_7),
    .io_out_bits_19_8(neuralNetsmidAndOutputWeightsMemory_io_out_bits_19_8),
    .io_out_bits_19_9(neuralNetsmidAndOutputWeightsMemory_io_out_bits_19_9),
    .io_out_bits_20_0(neuralNetsmidAndOutputWeightsMemory_io_out_bits_20_0),
    .io_out_bits_20_1(neuralNetsmidAndOutputWeightsMemory_io_out_bits_20_1),
    .io_out_bits_20_2(neuralNetsmidAndOutputWeightsMemory_io_out_bits_20_2),
    .io_out_bits_20_3(neuralNetsmidAndOutputWeightsMemory_io_out_bits_20_3),
    .io_out_bits_20_4(neuralNetsmidAndOutputWeightsMemory_io_out_bits_20_4),
    .io_out_bits_20_5(neuralNetsmidAndOutputWeightsMemory_io_out_bits_20_5),
    .io_out_bits_20_6(neuralNetsmidAndOutputWeightsMemory_io_out_bits_20_6),
    .io_out_bits_20_7(neuralNetsmidAndOutputWeightsMemory_io_out_bits_20_7),
    .io_out_bits_20_8(neuralNetsmidAndOutputWeightsMemory_io_out_bits_20_8),
    .io_out_bits_20_9(neuralNetsmidAndOutputWeightsMemory_io_out_bits_20_9)
  );
  MemoryBuffer_2 neuralNetsbiasVecsMemory ( // @[ConfigurationMemory.scala 84:40]
    .clock(neuralNetsbiasVecsMemory_clock),
    .reset(neuralNetsbiasVecsMemory_reset),
    .io_in_valid(neuralNetsbiasVecsMemory_io_in_valid),
    .io_in_bits(neuralNetsbiasVecsMemory_io_in_bits),
    .io_out_bits_0_0(neuralNetsbiasVecsMemory_io_out_bits_0_0),
    .io_out_bits_0_1(neuralNetsbiasVecsMemory_io_out_bits_0_1),
    .io_out_bits_0_2(neuralNetsbiasVecsMemory_io_out_bits_0_2),
    .io_out_bits_0_3(neuralNetsbiasVecsMemory_io_out_bits_0_3),
    .io_out_bits_0_4(neuralNetsbiasVecsMemory_io_out_bits_0_4),
    .io_out_bits_0_5(neuralNetsbiasVecsMemory_io_out_bits_0_5),
    .io_out_bits_0_6(neuralNetsbiasVecsMemory_io_out_bits_0_6),
    .io_out_bits_0_7(neuralNetsbiasVecsMemory_io_out_bits_0_7),
    .io_out_bits_0_8(neuralNetsbiasVecsMemory_io_out_bits_0_8),
    .io_out_bits_0_9(neuralNetsbiasVecsMemory_io_out_bits_0_9),
    .io_out_bits_1_0(neuralNetsbiasVecsMemory_io_out_bits_1_0),
    .io_out_bits_1_1(neuralNetsbiasVecsMemory_io_out_bits_1_1),
    .io_out_bits_1_2(neuralNetsbiasVecsMemory_io_out_bits_1_2),
    .io_out_bits_1_3(neuralNetsbiasVecsMemory_io_out_bits_1_3),
    .io_out_bits_1_4(neuralNetsbiasVecsMemory_io_out_bits_1_4),
    .io_out_bits_1_5(neuralNetsbiasVecsMemory_io_out_bits_1_5),
    .io_out_bits_1_6(neuralNetsbiasVecsMemory_io_out_bits_1_6),
    .io_out_bits_1_7(neuralNetsbiasVecsMemory_io_out_bits_1_7),
    .io_out_bits_1_8(neuralNetsbiasVecsMemory_io_out_bits_1_8),
    .io_out_bits_1_9(neuralNetsbiasVecsMemory_io_out_bits_1_9),
    .io_out_bits_2_0(neuralNetsbiasVecsMemory_io_out_bits_2_0),
    .io_out_bits_2_1(neuralNetsbiasVecsMemory_io_out_bits_2_1),
    .io_out_bits_2_2(neuralNetsbiasVecsMemory_io_out_bits_2_2),
    .io_out_bits_2_3(neuralNetsbiasVecsMemory_io_out_bits_2_3),
    .io_out_bits_2_4(neuralNetsbiasVecsMemory_io_out_bits_2_4),
    .io_out_bits_2_5(neuralNetsbiasVecsMemory_io_out_bits_2_5),
    .io_out_bits_2_6(neuralNetsbiasVecsMemory_io_out_bits_2_6),
    .io_out_bits_2_7(neuralNetsbiasVecsMemory_io_out_bits_2_7),
    .io_out_bits_2_8(neuralNetsbiasVecsMemory_io_out_bits_2_8),
    .io_out_bits_2_9(neuralNetsbiasVecsMemory_io_out_bits_2_9)
  );
  MemoryBuffer_3 neuralNetsoutputBiasMemory ( // @[ConfigurationMemory.scala 96:42]
    .clock(neuralNetsoutputBiasMemory_clock),
    .reset(neuralNetsoutputBiasMemory_reset),
    .io_in_valid(neuralNetsoutputBiasMemory_io_in_valid),
    .io_in_bits(neuralNetsoutputBiasMemory_io_in_bits),
    .io_out_bits_0_0(neuralNetsoutputBiasMemory_io_out_bits_0_0)
  );
  assign _T = io_in_bits_wraddr == 3'h0; // @[ConfigurationMemory.scala 64:68]
  assign _T_2 = io_in_bits_wraddr == 3'h1; // @[ConfigurationMemory.scala 76:75]
  assign _T_4 = io_in_bits_wraddr == 3'h2; // @[ConfigurationMemory.scala 87:64]
  assign _T_6 = io_in_bits_wraddr == 3'h3; // @[ConfigurationMemory.scala 99:66]
  assign _T_8 = io_in_bits_wraddr == 3'h4; // @[ConfigurationMemory.scala 105:29]
  assign _T_9 = io_in_valid & _T_8; // @[ConfigurationMemory.scala 105:20]
  assign _T_10 = $unsigned(io_in_bits_wrdata); // @[ConfigurationMemory.scala 105:90]
  assign _T_11 = _T_10[0]; // @[ConfigurationMemory.scala 105:92]
  assign io_out_bits_confneuralNetsinputWeights_0_0 = neuralNetsinputWeightsMemory_io_out_bits_0_0; // @[ConfigurationMemory.scala 65:42]
  assign io_out_bits_confneuralNetsinputWeights_0_1 = neuralNetsinputWeightsMemory_io_out_bits_0_1; // @[ConfigurationMemory.scala 65:42]
  assign io_out_bits_confneuralNetsinputWeights_0_2 = neuralNetsinputWeightsMemory_io_out_bits_0_2; // @[ConfigurationMemory.scala 65:42]
  assign io_out_bits_confneuralNetsinputWeights_0_3 = neuralNetsinputWeightsMemory_io_out_bits_0_3; // @[ConfigurationMemory.scala 65:42]
  assign io_out_bits_confneuralNetsinputWeights_1_0 = neuralNetsinputWeightsMemory_io_out_bits_1_0; // @[ConfigurationMemory.scala 65:42]
  assign io_out_bits_confneuralNetsinputWeights_1_1 = neuralNetsinputWeightsMemory_io_out_bits_1_1; // @[ConfigurationMemory.scala 65:42]
  assign io_out_bits_confneuralNetsinputWeights_1_2 = neuralNetsinputWeightsMemory_io_out_bits_1_2; // @[ConfigurationMemory.scala 65:42]
  assign io_out_bits_confneuralNetsinputWeights_1_3 = neuralNetsinputWeightsMemory_io_out_bits_1_3; // @[ConfigurationMemory.scala 65:42]
  assign io_out_bits_confneuralNetsinputWeights_2_0 = neuralNetsinputWeightsMemory_io_out_bits_2_0; // @[ConfigurationMemory.scala 65:42]
  assign io_out_bits_confneuralNetsinputWeights_2_1 = neuralNetsinputWeightsMemory_io_out_bits_2_1; // @[ConfigurationMemory.scala 65:42]
  assign io_out_bits_confneuralNetsinputWeights_2_2 = neuralNetsinputWeightsMemory_io_out_bits_2_2; // @[ConfigurationMemory.scala 65:42]
  assign io_out_bits_confneuralNetsinputWeights_2_3 = neuralNetsinputWeightsMemory_io_out_bits_2_3; // @[ConfigurationMemory.scala 65:42]
  assign io_out_bits_confneuralNetsinputWeights_3_0 = neuralNetsinputWeightsMemory_io_out_bits_3_0; // @[ConfigurationMemory.scala 65:42]
  assign io_out_bits_confneuralNetsinputWeights_3_1 = neuralNetsinputWeightsMemory_io_out_bits_3_1; // @[ConfigurationMemory.scala 65:42]
  assign io_out_bits_confneuralNetsinputWeights_3_2 = neuralNetsinputWeightsMemory_io_out_bits_3_2; // @[ConfigurationMemory.scala 65:42]
  assign io_out_bits_confneuralNetsinputWeights_3_3 = neuralNetsinputWeightsMemory_io_out_bits_3_3; // @[ConfigurationMemory.scala 65:42]
  assign io_out_bits_confneuralNetsinputWeights_4_0 = neuralNetsinputWeightsMemory_io_out_bits_4_0; // @[ConfigurationMemory.scala 65:42]
  assign io_out_bits_confneuralNetsinputWeights_4_1 = neuralNetsinputWeightsMemory_io_out_bits_4_1; // @[ConfigurationMemory.scala 65:42]
  assign io_out_bits_confneuralNetsinputWeights_4_2 = neuralNetsinputWeightsMemory_io_out_bits_4_2; // @[ConfigurationMemory.scala 65:42]
  assign io_out_bits_confneuralNetsinputWeights_4_3 = neuralNetsinputWeightsMemory_io_out_bits_4_3; // @[ConfigurationMemory.scala 65:42]
  assign io_out_bits_confneuralNetsinputWeights_5_0 = neuralNetsinputWeightsMemory_io_out_bits_5_0; // @[ConfigurationMemory.scala 65:42]
  assign io_out_bits_confneuralNetsinputWeights_5_1 = neuralNetsinputWeightsMemory_io_out_bits_5_1; // @[ConfigurationMemory.scala 65:42]
  assign io_out_bits_confneuralNetsinputWeights_5_2 = neuralNetsinputWeightsMemory_io_out_bits_5_2; // @[ConfigurationMemory.scala 65:42]
  assign io_out_bits_confneuralNetsinputWeights_5_3 = neuralNetsinputWeightsMemory_io_out_bits_5_3; // @[ConfigurationMemory.scala 65:42]
  assign io_out_bits_confneuralNetsinputWeights_6_0 = neuralNetsinputWeightsMemory_io_out_bits_6_0; // @[ConfigurationMemory.scala 65:42]
  assign io_out_bits_confneuralNetsinputWeights_6_1 = neuralNetsinputWeightsMemory_io_out_bits_6_1; // @[ConfigurationMemory.scala 65:42]
  assign io_out_bits_confneuralNetsinputWeights_6_2 = neuralNetsinputWeightsMemory_io_out_bits_6_2; // @[ConfigurationMemory.scala 65:42]
  assign io_out_bits_confneuralNetsinputWeights_6_3 = neuralNetsinputWeightsMemory_io_out_bits_6_3; // @[ConfigurationMemory.scala 65:42]
  assign io_out_bits_confneuralNetsinputWeights_7_0 = neuralNetsinputWeightsMemory_io_out_bits_7_0; // @[ConfigurationMemory.scala 65:42]
  assign io_out_bits_confneuralNetsinputWeights_7_1 = neuralNetsinputWeightsMemory_io_out_bits_7_1; // @[ConfigurationMemory.scala 65:42]
  assign io_out_bits_confneuralNetsinputWeights_7_2 = neuralNetsinputWeightsMemory_io_out_bits_7_2; // @[ConfigurationMemory.scala 65:42]
  assign io_out_bits_confneuralNetsinputWeights_7_3 = neuralNetsinputWeightsMemory_io_out_bits_7_3; // @[ConfigurationMemory.scala 65:42]
  assign io_out_bits_confneuralNetsinputWeights_8_0 = neuralNetsinputWeightsMemory_io_out_bits_8_0; // @[ConfigurationMemory.scala 65:42]
  assign io_out_bits_confneuralNetsinputWeights_8_1 = neuralNetsinputWeightsMemory_io_out_bits_8_1; // @[ConfigurationMemory.scala 65:42]
  assign io_out_bits_confneuralNetsinputWeights_8_2 = neuralNetsinputWeightsMemory_io_out_bits_8_2; // @[ConfigurationMemory.scala 65:42]
  assign io_out_bits_confneuralNetsinputWeights_8_3 = neuralNetsinputWeightsMemory_io_out_bits_8_3; // @[ConfigurationMemory.scala 65:42]
  assign io_out_bits_confneuralNetsinputWeights_9_0 = neuralNetsinputWeightsMemory_io_out_bits_9_0; // @[ConfigurationMemory.scala 65:42]
  assign io_out_bits_confneuralNetsinputWeights_9_1 = neuralNetsinputWeightsMemory_io_out_bits_9_1; // @[ConfigurationMemory.scala 65:42]
  assign io_out_bits_confneuralNetsinputWeights_9_2 = neuralNetsinputWeightsMemory_io_out_bits_9_2; // @[ConfigurationMemory.scala 65:42]
  assign io_out_bits_confneuralNetsinputWeights_9_3 = neuralNetsinputWeightsMemory_io_out_bits_9_3; // @[ConfigurationMemory.scala 65:42]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_0_0 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_0_0; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_0_1 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_0_1; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_0_2 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_0_2; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_0_3 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_0_3; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_0_4 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_0_4; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_0_5 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_0_5; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_0_6 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_0_6; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_0_7 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_0_7; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_0_8 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_0_8; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_0_9 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_0_9; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_1_0 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_1_0; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_1_1 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_1_1; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_1_2 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_1_2; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_1_3 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_1_3; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_1_4 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_1_4; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_1_5 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_1_5; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_1_6 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_1_6; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_1_7 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_1_7; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_1_8 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_1_8; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_1_9 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_1_9; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_2_0 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_2_0; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_2_1 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_2_1; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_2_2 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_2_2; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_2_3 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_2_3; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_2_4 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_2_4; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_2_5 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_2_5; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_2_6 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_2_6; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_2_7 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_2_7; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_2_8 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_2_8; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_2_9 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_2_9; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_3_0 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_3_0; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_3_1 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_3_1; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_3_2 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_3_2; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_3_3 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_3_3; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_3_4 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_3_4; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_3_5 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_3_5; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_3_6 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_3_6; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_3_7 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_3_7; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_3_8 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_3_8; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_3_9 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_3_9; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_4_0 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_4_0; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_4_1 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_4_1; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_4_2 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_4_2; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_4_3 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_4_3; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_4_4 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_4_4; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_4_5 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_4_5; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_4_6 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_4_6; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_4_7 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_4_7; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_4_8 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_4_8; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_4_9 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_4_9; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_5_0 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_5_0; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_5_1 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_5_1; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_5_2 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_5_2; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_5_3 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_5_3; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_5_4 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_5_4; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_5_5 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_5_5; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_5_6 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_5_6; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_5_7 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_5_7; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_5_8 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_5_8; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_5_9 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_5_9; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_6_0 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_6_0; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_6_1 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_6_1; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_6_2 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_6_2; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_6_3 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_6_3; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_6_4 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_6_4; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_6_5 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_6_5; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_6_6 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_6_6; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_6_7 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_6_7; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_6_8 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_6_8; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_6_9 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_6_9; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_7_0 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_7_0; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_7_1 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_7_1; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_7_2 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_7_2; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_7_3 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_7_3; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_7_4 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_7_4; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_7_5 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_7_5; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_7_6 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_7_6; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_7_7 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_7_7; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_7_8 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_7_8; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_7_9 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_7_9; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_8_0 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_8_0; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_8_1 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_8_1; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_8_2 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_8_2; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_8_3 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_8_3; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_8_4 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_8_4; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_8_5 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_8_5; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_8_6 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_8_6; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_8_7 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_8_7; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_8_8 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_8_8; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_8_9 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_8_9; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_9_0 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_9_0; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_9_1 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_9_1; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_9_2 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_9_2; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_9_3 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_9_3; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_9_4 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_9_4; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_9_5 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_9_5; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_9_6 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_9_6; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_9_7 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_9_7; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_9_8 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_9_8; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_9_9 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_9_9; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_10_0 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_10_0; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_10_1 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_10_1; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_10_2 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_10_2; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_10_3 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_10_3; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_10_4 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_10_4; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_10_5 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_10_5; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_10_6 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_10_6; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_10_7 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_10_7; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_10_8 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_10_8; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_10_9 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_10_9; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_11_0 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_11_0; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_11_1 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_11_1; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_11_2 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_11_2; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_11_3 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_11_3; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_11_4 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_11_4; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_11_5 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_11_5; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_11_6 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_11_6; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_11_7 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_11_7; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_11_8 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_11_8; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_11_9 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_11_9; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_12_0 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_12_0; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_12_1 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_12_1; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_12_2 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_12_2; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_12_3 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_12_3; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_12_4 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_12_4; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_12_5 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_12_5; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_12_6 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_12_6; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_12_7 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_12_7; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_12_8 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_12_8; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_12_9 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_12_9; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_13_0 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_13_0; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_13_1 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_13_1; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_13_2 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_13_2; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_13_3 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_13_3; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_13_4 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_13_4; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_13_5 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_13_5; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_13_6 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_13_6; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_13_7 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_13_7; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_13_8 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_13_8; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_13_9 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_13_9; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_14_0 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_14_0; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_14_1 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_14_1; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_14_2 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_14_2; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_14_3 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_14_3; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_14_4 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_14_4; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_14_5 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_14_5; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_14_6 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_14_6; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_14_7 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_14_7; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_14_8 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_14_8; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_14_9 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_14_9; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_15_0 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_15_0; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_15_1 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_15_1; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_15_2 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_15_2; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_15_3 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_15_3; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_15_4 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_15_4; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_15_5 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_15_5; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_15_6 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_15_6; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_15_7 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_15_7; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_15_8 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_15_8; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_15_9 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_15_9; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_16_0 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_16_0; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_16_1 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_16_1; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_16_2 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_16_2; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_16_3 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_16_3; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_16_4 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_16_4; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_16_5 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_16_5; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_16_6 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_16_6; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_16_7 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_16_7; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_16_8 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_16_8; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_16_9 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_16_9; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_17_0 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_17_0; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_17_1 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_17_1; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_17_2 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_17_2; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_17_3 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_17_3; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_17_4 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_17_4; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_17_5 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_17_5; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_17_6 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_17_6; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_17_7 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_17_7; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_17_8 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_17_8; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_17_9 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_17_9; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_18_0 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_18_0; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_18_1 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_18_1; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_18_2 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_18_2; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_18_3 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_18_3; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_18_4 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_18_4; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_18_5 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_18_5; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_18_6 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_18_6; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_18_7 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_18_7; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_18_8 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_18_8; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_18_9 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_18_9; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_19_0 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_19_0; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_19_1 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_19_1; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_19_2 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_19_2; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_19_3 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_19_3; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_19_4 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_19_4; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_19_5 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_19_5; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_19_6 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_19_6; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_19_7 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_19_7; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_19_8 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_19_8; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_19_9 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_19_9; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_20_0 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_20_0; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_20_1 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_20_1; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_20_2 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_20_2; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_20_3 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_20_3; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_20_4 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_20_4; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_20_5 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_20_5; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_20_6 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_20_6; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_20_7 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_20_7; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_20_8 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_20_8; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsmidAndOutputWeights_20_9 = neuralNetsmidAndOutputWeightsMemory_io_out_bits_20_9; // @[ConfigurationMemory.scala 77:49]
  assign io_out_bits_confneuralNetsbiasVecs_0_0 = neuralNetsbiasVecsMemory_io_out_bits_0_0; // @[ConfigurationMemory.scala 88:38]
  assign io_out_bits_confneuralNetsbiasVecs_0_1 = neuralNetsbiasVecsMemory_io_out_bits_0_1; // @[ConfigurationMemory.scala 88:38]
  assign io_out_bits_confneuralNetsbiasVecs_0_2 = neuralNetsbiasVecsMemory_io_out_bits_0_2; // @[ConfigurationMemory.scala 88:38]
  assign io_out_bits_confneuralNetsbiasVecs_0_3 = neuralNetsbiasVecsMemory_io_out_bits_0_3; // @[ConfigurationMemory.scala 88:38]
  assign io_out_bits_confneuralNetsbiasVecs_0_4 = neuralNetsbiasVecsMemory_io_out_bits_0_4; // @[ConfigurationMemory.scala 88:38]
  assign io_out_bits_confneuralNetsbiasVecs_0_5 = neuralNetsbiasVecsMemory_io_out_bits_0_5; // @[ConfigurationMemory.scala 88:38]
  assign io_out_bits_confneuralNetsbiasVecs_0_6 = neuralNetsbiasVecsMemory_io_out_bits_0_6; // @[ConfigurationMemory.scala 88:38]
  assign io_out_bits_confneuralNetsbiasVecs_0_7 = neuralNetsbiasVecsMemory_io_out_bits_0_7; // @[ConfigurationMemory.scala 88:38]
  assign io_out_bits_confneuralNetsbiasVecs_0_8 = neuralNetsbiasVecsMemory_io_out_bits_0_8; // @[ConfigurationMemory.scala 88:38]
  assign io_out_bits_confneuralNetsbiasVecs_0_9 = neuralNetsbiasVecsMemory_io_out_bits_0_9; // @[ConfigurationMemory.scala 88:38]
  assign io_out_bits_confneuralNetsbiasVecs_1_0 = neuralNetsbiasVecsMemory_io_out_bits_1_0; // @[ConfigurationMemory.scala 88:38]
  assign io_out_bits_confneuralNetsbiasVecs_1_1 = neuralNetsbiasVecsMemory_io_out_bits_1_1; // @[ConfigurationMemory.scala 88:38]
  assign io_out_bits_confneuralNetsbiasVecs_1_2 = neuralNetsbiasVecsMemory_io_out_bits_1_2; // @[ConfigurationMemory.scala 88:38]
  assign io_out_bits_confneuralNetsbiasVecs_1_3 = neuralNetsbiasVecsMemory_io_out_bits_1_3; // @[ConfigurationMemory.scala 88:38]
  assign io_out_bits_confneuralNetsbiasVecs_1_4 = neuralNetsbiasVecsMemory_io_out_bits_1_4; // @[ConfigurationMemory.scala 88:38]
  assign io_out_bits_confneuralNetsbiasVecs_1_5 = neuralNetsbiasVecsMemory_io_out_bits_1_5; // @[ConfigurationMemory.scala 88:38]
  assign io_out_bits_confneuralNetsbiasVecs_1_6 = neuralNetsbiasVecsMemory_io_out_bits_1_6; // @[ConfigurationMemory.scala 88:38]
  assign io_out_bits_confneuralNetsbiasVecs_1_7 = neuralNetsbiasVecsMemory_io_out_bits_1_7; // @[ConfigurationMemory.scala 88:38]
  assign io_out_bits_confneuralNetsbiasVecs_1_8 = neuralNetsbiasVecsMemory_io_out_bits_1_8; // @[ConfigurationMemory.scala 88:38]
  assign io_out_bits_confneuralNetsbiasVecs_1_9 = neuralNetsbiasVecsMemory_io_out_bits_1_9; // @[ConfigurationMemory.scala 88:38]
  assign io_out_bits_confneuralNetsbiasVecs_2_0 = neuralNetsbiasVecsMemory_io_out_bits_2_0; // @[ConfigurationMemory.scala 88:38]
  assign io_out_bits_confneuralNetsbiasVecs_2_1 = neuralNetsbiasVecsMemory_io_out_bits_2_1; // @[ConfigurationMemory.scala 88:38]
  assign io_out_bits_confneuralNetsbiasVecs_2_2 = neuralNetsbiasVecsMemory_io_out_bits_2_2; // @[ConfigurationMemory.scala 88:38]
  assign io_out_bits_confneuralNetsbiasVecs_2_3 = neuralNetsbiasVecsMemory_io_out_bits_2_3; // @[ConfigurationMemory.scala 88:38]
  assign io_out_bits_confneuralNetsbiasVecs_2_4 = neuralNetsbiasVecsMemory_io_out_bits_2_4; // @[ConfigurationMemory.scala 88:38]
  assign io_out_bits_confneuralNetsbiasVecs_2_5 = neuralNetsbiasVecsMemory_io_out_bits_2_5; // @[ConfigurationMemory.scala 88:38]
  assign io_out_bits_confneuralNetsbiasVecs_2_6 = neuralNetsbiasVecsMemory_io_out_bits_2_6; // @[ConfigurationMemory.scala 88:38]
  assign io_out_bits_confneuralNetsbiasVecs_2_7 = neuralNetsbiasVecsMemory_io_out_bits_2_7; // @[ConfigurationMemory.scala 88:38]
  assign io_out_bits_confneuralNetsbiasVecs_2_8 = neuralNetsbiasVecsMemory_io_out_bits_2_8; // @[ConfigurationMemory.scala 88:38]
  assign io_out_bits_confneuralNetsbiasVecs_2_9 = neuralNetsbiasVecsMemory_io_out_bits_2_9; // @[ConfigurationMemory.scala 88:38]
  assign io_out_bits_confneuralNetsoutputBias_0 = neuralNetsoutputBiasMemory_io_out_bits_0_0; // @[ConfigurationMemory.scala 100:40]
  assign io_out_bits_confInputMuxSel = inputMuxSel; // @[ConfigurationMemory.scala 106:31]
  assign neuralNetsinputWeightsMemory_clock = clock;
  assign neuralNetsinputWeightsMemory_reset = reset;
  assign neuralNetsinputWeightsMemory_io_in_valid = io_in_valid & _T; // @[ConfigurationMemory.scala 64:44]
  assign neuralNetsinputWeightsMemory_io_in_bits = io_in_bits_wrdata; // @[ConfigurationMemory.scala 62:43]
  assign neuralNetsmidAndOutputWeightsMemory_clock = clock;
  assign neuralNetsmidAndOutputWeightsMemory_reset = reset;
  assign neuralNetsmidAndOutputWeightsMemory_io_in_valid = io_in_valid & _T_2; // @[ConfigurationMemory.scala 76:51]
  assign neuralNetsmidAndOutputWeightsMemory_io_in_bits = io_in_bits_wrdata; // @[ConfigurationMemory.scala 74:50]
  assign neuralNetsbiasVecsMemory_clock = clock;
  assign neuralNetsbiasVecsMemory_reset = reset;
  assign neuralNetsbiasVecsMemory_io_in_valid = io_in_valid & _T_4; // @[ConfigurationMemory.scala 87:40]
  assign neuralNetsbiasVecsMemory_io_in_bits = io_in_bits_wrdata; // @[ConfigurationMemory.scala 85:39]
  assign neuralNetsoutputBiasMemory_clock = clock;
  assign neuralNetsoutputBiasMemory_reset = reset;
  assign neuralNetsoutputBiasMemory_io_in_valid = io_in_valid & _T_6; // @[ConfigurationMemory.scala 99:42]
  assign neuralNetsoutputBiasMemory_io_in_bits = io_in_bits_wrdata; // @[ConfigurationMemory.scala 97:41]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  inputMuxSel = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      inputMuxSel <= 1'h0;
    end else begin
      if (_T_9) begin
        inputMuxSel <= _T_11;
      end
    end
  end
endmodule
module TLWellnessDataPathBlock(
  input         clock,
  input         reset,
  output        in_ready,
  input         in_valid,
  input  [63:0] in_bits_data,
  input         in_bits_last,
  input         out_ready,
  output        out_valid,
  output [63:0] out_bits_data,
  output        out_bits_last,
  output        in2_ready,
  input         in2_valid,
  input  [63:0] in2_bits_data,
  input         in2_bits_last,
  input         streamIn_valid,
  input  [31:0] streamIn_bits,
  input         streamIn_sync
);
  wire  converter_auto_in_ready; // @[Nodes.scala 106:31]
  wire  converter_auto_in_valid; // @[Nodes.scala 106:31]
  wire [63:0] converter_auto_in_bits_data; // @[Nodes.scala 106:31]
  wire  converter_auto_in_bits_last; // @[Nodes.scala 106:31]
  wire  converter_auto_out_ready; // @[Nodes.scala 106:31]
  wire  converter_auto_out_valid; // @[Nodes.scala 106:31]
  wire [63:0] converter_auto_out_bits_data; // @[Nodes.scala 106:31]
  wire  converter_auto_out_bits_last; // @[Nodes.scala 106:31]
  wire  converter_1_auto_in_ready; // @[Nodes.scala 142:31]
  wire  converter_1_auto_in_valid; // @[Nodes.scala 142:31]
  wire [63:0] converter_1_auto_in_bits_data; // @[Nodes.scala 142:31]
  wire  converter_1_auto_in_bits_last; // @[Nodes.scala 142:31]
  wire  converter_1_auto_out_ready; // @[Nodes.scala 142:31]
  wire  converter_1_auto_out_valid; // @[Nodes.scala 142:31]
  wire [63:0] converter_1_auto_out_bits_data; // @[Nodes.scala 142:31]
  wire  converter_1_auto_out_bits_last; // @[Nodes.scala 142:31]
  wire  converter_2_auto_in_ready; // @[Nodes.scala 142:31]
  wire  converter_2_auto_in_valid; // @[Nodes.scala 142:31]
  wire [63:0] converter_2_auto_in_bits_data; // @[Nodes.scala 142:31]
  wire  converter_2_auto_in_bits_last; // @[Nodes.scala 142:31]
  wire  converter_2_auto_out_ready; // @[Nodes.scala 142:31]
  wire  converter_2_auto_out_valid; // @[Nodes.scala 142:31]
  wire [63:0] converter_2_auto_out_bits_data; // @[Nodes.scala 142:31]
  wire  converter_2_auto_out_bits_last; // @[Nodes.scala 142:31]
  wire  wellness_clock; // @[Wellness.scala 388:26]
  wire  wellness_reset; // @[Wellness.scala 388:26]
  wire  wellness_io_streamIn_valid; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_streamIn_bits; // @[Wellness.scala 388:26]
  wire  wellness_io_in_valid; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_in_bits; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsinputWeights_0_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsinputWeights_0_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsinputWeights_0_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsinputWeights_0_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsinputWeights_1_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsinputWeights_1_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsinputWeights_1_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsinputWeights_1_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsinputWeights_2_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsinputWeights_2_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsinputWeights_2_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsinputWeights_2_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsinputWeights_3_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsinputWeights_3_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsinputWeights_3_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsinputWeights_3_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsinputWeights_4_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsinputWeights_4_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsinputWeights_4_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsinputWeights_4_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsinputWeights_5_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsinputWeights_5_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsinputWeights_5_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsinputWeights_5_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsinputWeights_6_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsinputWeights_6_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsinputWeights_6_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsinputWeights_6_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsinputWeights_7_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsinputWeights_7_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsinputWeights_7_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsinputWeights_7_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsinputWeights_8_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsinputWeights_8_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsinputWeights_8_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsinputWeights_8_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsinputWeights_9_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsinputWeights_9_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsinputWeights_9_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsinputWeights_9_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_0_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_0_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_0_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_0_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_0_4; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_0_5; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_0_6; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_0_7; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_0_8; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_0_9; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_1_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_1_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_1_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_1_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_1_4; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_1_5; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_1_6; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_1_7; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_1_8; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_1_9; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_2_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_2_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_2_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_2_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_2_4; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_2_5; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_2_6; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_2_7; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_2_8; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_2_9; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_3_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_3_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_3_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_3_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_3_4; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_3_5; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_3_6; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_3_7; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_3_8; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_3_9; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_4_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_4_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_4_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_4_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_4_4; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_4_5; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_4_6; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_4_7; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_4_8; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_4_9; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_5_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_5_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_5_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_5_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_5_4; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_5_5; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_5_6; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_5_7; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_5_8; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_5_9; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_6_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_6_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_6_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_6_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_6_4; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_6_5; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_6_6; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_6_7; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_6_8; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_6_9; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_7_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_7_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_7_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_7_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_7_4; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_7_5; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_7_6; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_7_7; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_7_8; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_7_9; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_8_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_8_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_8_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_8_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_8_4; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_8_5; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_8_6; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_8_7; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_8_8; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_8_9; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_9_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_9_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_9_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_9_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_9_4; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_9_5; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_9_6; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_9_7; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_9_8; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_9_9; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_10_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_10_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_10_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_10_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_10_4; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_10_5; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_10_6; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_10_7; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_10_8; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_10_9; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_11_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_11_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_11_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_11_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_11_4; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_11_5; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_11_6; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_11_7; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_11_8; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_11_9; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_12_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_12_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_12_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_12_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_12_4; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_12_5; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_12_6; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_12_7; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_12_8; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_12_9; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_13_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_13_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_13_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_13_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_13_4; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_13_5; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_13_6; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_13_7; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_13_8; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_13_9; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_14_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_14_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_14_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_14_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_14_4; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_14_5; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_14_6; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_14_7; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_14_8; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_14_9; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_15_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_15_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_15_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_15_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_15_4; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_15_5; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_15_6; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_15_7; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_15_8; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_15_9; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_16_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_16_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_16_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_16_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_16_4; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_16_5; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_16_6; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_16_7; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_16_8; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_16_9; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_17_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_17_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_17_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_17_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_17_4; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_17_5; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_17_6; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_17_7; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_17_8; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_17_9; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_18_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_18_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_18_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_18_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_18_4; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_18_5; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_18_6; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_18_7; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_18_8; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_18_9; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_19_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_19_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_19_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_19_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_19_4; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_19_5; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_19_6; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_19_7; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_19_8; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_19_9; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_20_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_20_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_20_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_20_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_20_4; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_20_5; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_20_6; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_20_7; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_20_8; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_20_9; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVecs_0_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVecs_0_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVecs_0_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVecs_0_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVecs_0_4; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVecs_0_5; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVecs_0_6; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVecs_0_7; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVecs_0_8; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVecs_0_9; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVecs_1_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVecs_1_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVecs_1_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVecs_1_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVecs_1_4; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVecs_1_5; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVecs_1_6; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVecs_1_7; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVecs_1_8; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVecs_1_9; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVecs_2_0; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVecs_2_1; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVecs_2_2; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVecs_2_3; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVecs_2_4; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVecs_2_5; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVecs_2_6; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVecs_2_7; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVecs_2_8; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsbiasVecs_2_9; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_inConf_bits_confneuralNetsoutputBias_0; // @[Wellness.scala 388:26]
  wire  wellness_io_inConf_bits_confInputMuxSel; // @[Wellness.scala 388:26]
  wire  wellness_io_out_valid; // @[Wellness.scala 388:26]
  wire  wellness_io_out_bits; // @[Wellness.scala 388:26]
  wire [31:0] wellness_io_rawVotes; // @[Wellness.scala 388:26]
  wire  configurationMemory_clock; // @[Wellness.scala 398:37]
  wire  configurationMemory_reset; // @[Wellness.scala 398:37]
  wire  configurationMemory_io_in_valid; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_in_bits_wrdata; // @[Wellness.scala 398:37]
  wire [2:0] configurationMemory_io_in_bits_wraddr; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsinputWeights_0_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsinputWeights_0_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsinputWeights_0_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsinputWeights_0_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsinputWeights_1_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsinputWeights_1_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsinputWeights_1_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsinputWeights_1_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsinputWeights_2_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsinputWeights_2_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsinputWeights_2_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsinputWeights_2_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsinputWeights_3_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsinputWeights_3_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsinputWeights_3_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsinputWeights_3_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsinputWeights_4_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsinputWeights_4_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsinputWeights_4_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsinputWeights_4_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsinputWeights_5_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsinputWeights_5_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsinputWeights_5_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsinputWeights_5_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsinputWeights_6_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsinputWeights_6_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsinputWeights_6_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsinputWeights_6_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsinputWeights_7_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsinputWeights_7_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsinputWeights_7_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsinputWeights_7_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsinputWeights_8_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsinputWeights_8_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsinputWeights_8_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsinputWeights_8_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsinputWeights_9_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsinputWeights_9_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsinputWeights_9_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsinputWeights_9_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_0_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_0_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_0_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_0_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_0_4; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_0_5; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_0_6; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_0_7; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_0_8; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_0_9; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_1_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_1_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_1_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_1_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_1_4; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_1_5; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_1_6; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_1_7; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_1_8; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_1_9; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_2_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_2_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_2_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_2_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_2_4; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_2_5; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_2_6; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_2_7; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_2_8; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_2_9; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_3_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_3_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_3_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_3_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_3_4; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_3_5; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_3_6; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_3_7; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_3_8; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_3_9; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_4_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_4_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_4_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_4_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_4_4; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_4_5; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_4_6; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_4_7; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_4_8; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_4_9; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_5_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_5_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_5_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_5_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_5_4; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_5_5; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_5_6; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_5_7; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_5_8; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_5_9; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_6_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_6_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_6_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_6_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_6_4; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_6_5; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_6_6; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_6_7; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_6_8; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_6_9; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_7_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_7_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_7_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_7_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_7_4; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_7_5; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_7_6; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_7_7; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_7_8; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_7_9; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_8_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_8_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_8_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_8_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_8_4; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_8_5; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_8_6; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_8_7; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_8_8; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_8_9; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_9_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_9_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_9_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_9_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_9_4; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_9_5; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_9_6; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_9_7; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_9_8; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_9_9; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_10_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_10_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_10_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_10_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_10_4; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_10_5; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_10_6; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_10_7; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_10_8; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_10_9; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_11_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_11_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_11_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_11_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_11_4; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_11_5; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_11_6; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_11_7; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_11_8; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_11_9; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_12_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_12_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_12_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_12_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_12_4; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_12_5; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_12_6; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_12_7; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_12_8; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_12_9; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_13_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_13_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_13_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_13_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_13_4; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_13_5; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_13_6; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_13_7; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_13_8; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_13_9; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_14_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_14_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_14_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_14_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_14_4; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_14_5; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_14_6; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_14_7; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_14_8; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_14_9; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_15_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_15_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_15_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_15_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_15_4; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_15_5; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_15_6; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_15_7; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_15_8; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_15_9; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_16_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_16_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_16_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_16_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_16_4; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_16_5; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_16_6; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_16_7; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_16_8; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_16_9; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_17_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_17_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_17_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_17_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_17_4; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_17_5; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_17_6; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_17_7; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_17_8; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_17_9; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_18_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_18_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_18_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_18_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_18_4; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_18_5; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_18_6; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_18_7; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_18_8; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_18_9; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_19_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_19_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_19_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_19_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_19_4; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_19_5; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_19_6; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_19_7; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_19_8; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_19_9; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_20_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_20_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_20_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_20_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_20_4; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_20_5; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_20_6; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_20_7; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_20_8; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_20_9; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVecs_0_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVecs_0_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVecs_0_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVecs_0_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVecs_0_4; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVecs_0_5; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVecs_0_6; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVecs_0_7; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVecs_0_8; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVecs_0_9; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVecs_1_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVecs_1_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVecs_1_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVecs_1_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVecs_1_4; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVecs_1_5; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVecs_1_6; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVecs_1_7; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVecs_1_8; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVecs_1_9; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVecs_2_0; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVecs_2_1; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVecs_2_2; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVecs_2_3; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVecs_2_4; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVecs_2_5; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVecs_2_6; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVecs_2_7; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVecs_2_8; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsbiasVecs_2_9; // @[Wellness.scala 398:37]
  wire [31:0] configurationMemory_io_out_bits_confneuralNetsoutputBias_0; // @[Wellness.scala 398:37]
  wire  configurationMemory_io_out_bits_confInputMuxSel; // @[Wellness.scala 398:37]
  wire [63:0] in_1_bits_data; // @[Nodes.scala 333:76 LazyModule.scala 167:31]
  wire [63:0] _T_4; // @[Wellness.scala 408:49]
  wire [31:0] _T_5; // @[Wellness.scala 411:83]
  wire [32:0] _T_6; // @[Cat.scala 30:58]
  wire [63:0] inConf_bits_data; // @[Nodes.scala 333:76 LazyModule.scala 167:31]
  wire [31:0] _T_7; // @[Wellness.scala 418:62]
  wire [31:0] _GEN_0; // @[Wellness.scala 408:49 Wellness.scala 408:49]
  AXI4StreamToBundleBridge converter ( // @[Nodes.scala 106:31]
    .auto_in_ready(converter_auto_in_ready),
    .auto_in_valid(converter_auto_in_valid),
    .auto_in_bits_data(converter_auto_in_bits_data),
    .auto_in_bits_last(converter_auto_in_bits_last),
    .auto_out_ready(converter_auto_out_ready),
    .auto_out_valid(converter_auto_out_valid),
    .auto_out_bits_data(converter_auto_out_bits_data),
    .auto_out_bits_last(converter_auto_out_bits_last)
  );
  AXI4StreamToBundleBridge converter_1 ( // @[Nodes.scala 142:31]
    .auto_in_ready(converter_1_auto_in_ready),
    .auto_in_valid(converter_1_auto_in_valid),
    .auto_in_bits_data(converter_1_auto_in_bits_data),
    .auto_in_bits_last(converter_1_auto_in_bits_last),
    .auto_out_ready(converter_1_auto_out_ready),
    .auto_out_valid(converter_1_auto_out_valid),
    .auto_out_bits_data(converter_1_auto_out_bits_data),
    .auto_out_bits_last(converter_1_auto_out_bits_last)
  );
  AXI4StreamToBundleBridge converter_2 ( // @[Nodes.scala 142:31]
    .auto_in_ready(converter_2_auto_in_ready),
    .auto_in_valid(converter_2_auto_in_valid),
    .auto_in_bits_data(converter_2_auto_in_bits_data),
    .auto_in_bits_last(converter_2_auto_in_bits_last),
    .auto_out_ready(converter_2_auto_out_ready),
    .auto_out_valid(converter_2_auto_out_valid),
    .auto_out_bits_data(converter_2_auto_out_bits_data),
    .auto_out_bits_last(converter_2_auto_out_bits_last)
  );
  WellnessModule wellness ( // @[Wellness.scala 388:26]
    .clock(wellness_clock),
    .reset(wellness_reset),
    .io_streamIn_valid(wellness_io_streamIn_valid),
    .io_streamIn_bits(wellness_io_streamIn_bits),
    .io_in_valid(wellness_io_in_valid),
    .io_in_bits(wellness_io_in_bits),
    .io_inConf_bits_confneuralNetsinputWeights_0_0(wellness_io_inConf_bits_confneuralNetsinputWeights_0_0),
    .io_inConf_bits_confneuralNetsinputWeights_0_1(wellness_io_inConf_bits_confneuralNetsinputWeights_0_1),
    .io_inConf_bits_confneuralNetsinputWeights_0_2(wellness_io_inConf_bits_confneuralNetsinputWeights_0_2),
    .io_inConf_bits_confneuralNetsinputWeights_0_3(wellness_io_inConf_bits_confneuralNetsinputWeights_0_3),
    .io_inConf_bits_confneuralNetsinputWeights_1_0(wellness_io_inConf_bits_confneuralNetsinputWeights_1_0),
    .io_inConf_bits_confneuralNetsinputWeights_1_1(wellness_io_inConf_bits_confneuralNetsinputWeights_1_1),
    .io_inConf_bits_confneuralNetsinputWeights_1_2(wellness_io_inConf_bits_confneuralNetsinputWeights_1_2),
    .io_inConf_bits_confneuralNetsinputWeights_1_3(wellness_io_inConf_bits_confneuralNetsinputWeights_1_3),
    .io_inConf_bits_confneuralNetsinputWeights_2_0(wellness_io_inConf_bits_confneuralNetsinputWeights_2_0),
    .io_inConf_bits_confneuralNetsinputWeights_2_1(wellness_io_inConf_bits_confneuralNetsinputWeights_2_1),
    .io_inConf_bits_confneuralNetsinputWeights_2_2(wellness_io_inConf_bits_confneuralNetsinputWeights_2_2),
    .io_inConf_bits_confneuralNetsinputWeights_2_3(wellness_io_inConf_bits_confneuralNetsinputWeights_2_3),
    .io_inConf_bits_confneuralNetsinputWeights_3_0(wellness_io_inConf_bits_confneuralNetsinputWeights_3_0),
    .io_inConf_bits_confneuralNetsinputWeights_3_1(wellness_io_inConf_bits_confneuralNetsinputWeights_3_1),
    .io_inConf_bits_confneuralNetsinputWeights_3_2(wellness_io_inConf_bits_confneuralNetsinputWeights_3_2),
    .io_inConf_bits_confneuralNetsinputWeights_3_3(wellness_io_inConf_bits_confneuralNetsinputWeights_3_3),
    .io_inConf_bits_confneuralNetsinputWeights_4_0(wellness_io_inConf_bits_confneuralNetsinputWeights_4_0),
    .io_inConf_bits_confneuralNetsinputWeights_4_1(wellness_io_inConf_bits_confneuralNetsinputWeights_4_1),
    .io_inConf_bits_confneuralNetsinputWeights_4_2(wellness_io_inConf_bits_confneuralNetsinputWeights_4_2),
    .io_inConf_bits_confneuralNetsinputWeights_4_3(wellness_io_inConf_bits_confneuralNetsinputWeights_4_3),
    .io_inConf_bits_confneuralNetsinputWeights_5_0(wellness_io_inConf_bits_confneuralNetsinputWeights_5_0),
    .io_inConf_bits_confneuralNetsinputWeights_5_1(wellness_io_inConf_bits_confneuralNetsinputWeights_5_1),
    .io_inConf_bits_confneuralNetsinputWeights_5_2(wellness_io_inConf_bits_confneuralNetsinputWeights_5_2),
    .io_inConf_bits_confneuralNetsinputWeights_5_3(wellness_io_inConf_bits_confneuralNetsinputWeights_5_3),
    .io_inConf_bits_confneuralNetsinputWeights_6_0(wellness_io_inConf_bits_confneuralNetsinputWeights_6_0),
    .io_inConf_bits_confneuralNetsinputWeights_6_1(wellness_io_inConf_bits_confneuralNetsinputWeights_6_1),
    .io_inConf_bits_confneuralNetsinputWeights_6_2(wellness_io_inConf_bits_confneuralNetsinputWeights_6_2),
    .io_inConf_bits_confneuralNetsinputWeights_6_3(wellness_io_inConf_bits_confneuralNetsinputWeights_6_3),
    .io_inConf_bits_confneuralNetsinputWeights_7_0(wellness_io_inConf_bits_confneuralNetsinputWeights_7_0),
    .io_inConf_bits_confneuralNetsinputWeights_7_1(wellness_io_inConf_bits_confneuralNetsinputWeights_7_1),
    .io_inConf_bits_confneuralNetsinputWeights_7_2(wellness_io_inConf_bits_confneuralNetsinputWeights_7_2),
    .io_inConf_bits_confneuralNetsinputWeights_7_3(wellness_io_inConf_bits_confneuralNetsinputWeights_7_3),
    .io_inConf_bits_confneuralNetsinputWeights_8_0(wellness_io_inConf_bits_confneuralNetsinputWeights_8_0),
    .io_inConf_bits_confneuralNetsinputWeights_8_1(wellness_io_inConf_bits_confneuralNetsinputWeights_8_1),
    .io_inConf_bits_confneuralNetsinputWeights_8_2(wellness_io_inConf_bits_confneuralNetsinputWeights_8_2),
    .io_inConf_bits_confneuralNetsinputWeights_8_3(wellness_io_inConf_bits_confneuralNetsinputWeights_8_3),
    .io_inConf_bits_confneuralNetsinputWeights_9_0(wellness_io_inConf_bits_confneuralNetsinputWeights_9_0),
    .io_inConf_bits_confneuralNetsinputWeights_9_1(wellness_io_inConf_bits_confneuralNetsinputWeights_9_1),
    .io_inConf_bits_confneuralNetsinputWeights_9_2(wellness_io_inConf_bits_confneuralNetsinputWeights_9_2),
    .io_inConf_bits_confneuralNetsinputWeights_9_3(wellness_io_inConf_bits_confneuralNetsinputWeights_9_3),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_0_0(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_0_0),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_0_1(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_0_1),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_0_2(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_0_2),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_0_3(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_0_3),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_0_4(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_0_4),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_0_5(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_0_5),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_0_6(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_0_6),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_0_7(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_0_7),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_0_8(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_0_8),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_0_9(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_0_9),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_1_0(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_1_0),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_1_1(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_1_1),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_1_2(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_1_2),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_1_3(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_1_3),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_1_4(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_1_4),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_1_5(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_1_5),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_1_6(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_1_6),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_1_7(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_1_7),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_1_8(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_1_8),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_1_9(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_1_9),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_2_0(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_2_0),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_2_1(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_2_1),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_2_2(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_2_2),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_2_3(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_2_3),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_2_4(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_2_4),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_2_5(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_2_5),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_2_6(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_2_6),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_2_7(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_2_7),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_2_8(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_2_8),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_2_9(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_2_9),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_3_0(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_3_0),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_3_1(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_3_1),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_3_2(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_3_2),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_3_3(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_3_3),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_3_4(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_3_4),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_3_5(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_3_5),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_3_6(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_3_6),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_3_7(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_3_7),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_3_8(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_3_8),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_3_9(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_3_9),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_4_0(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_4_0),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_4_1(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_4_1),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_4_2(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_4_2),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_4_3(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_4_3),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_4_4(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_4_4),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_4_5(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_4_5),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_4_6(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_4_6),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_4_7(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_4_7),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_4_8(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_4_8),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_4_9(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_4_9),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_5_0(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_5_0),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_5_1(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_5_1),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_5_2(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_5_2),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_5_3(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_5_3),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_5_4(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_5_4),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_5_5(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_5_5),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_5_6(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_5_6),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_5_7(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_5_7),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_5_8(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_5_8),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_5_9(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_5_9),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_6_0(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_6_0),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_6_1(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_6_1),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_6_2(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_6_2),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_6_3(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_6_3),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_6_4(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_6_4),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_6_5(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_6_5),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_6_6(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_6_6),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_6_7(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_6_7),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_6_8(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_6_8),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_6_9(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_6_9),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_7_0(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_7_0),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_7_1(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_7_1),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_7_2(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_7_2),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_7_3(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_7_3),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_7_4(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_7_4),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_7_5(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_7_5),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_7_6(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_7_6),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_7_7(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_7_7),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_7_8(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_7_8),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_7_9(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_7_9),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_8_0(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_8_0),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_8_1(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_8_1),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_8_2(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_8_2),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_8_3(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_8_3),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_8_4(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_8_4),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_8_5(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_8_5),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_8_6(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_8_6),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_8_7(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_8_7),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_8_8(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_8_8),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_8_9(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_8_9),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_9_0(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_9_0),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_9_1(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_9_1),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_9_2(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_9_2),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_9_3(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_9_3),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_9_4(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_9_4),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_9_5(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_9_5),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_9_6(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_9_6),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_9_7(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_9_7),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_9_8(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_9_8),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_9_9(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_9_9),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_10_0(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_10_0),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_10_1(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_10_1),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_10_2(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_10_2),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_10_3(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_10_3),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_10_4(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_10_4),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_10_5(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_10_5),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_10_6(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_10_6),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_10_7(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_10_7),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_10_8(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_10_8),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_10_9(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_10_9),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_11_0(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_11_0),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_11_1(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_11_1),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_11_2(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_11_2),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_11_3(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_11_3),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_11_4(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_11_4),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_11_5(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_11_5),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_11_6(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_11_6),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_11_7(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_11_7),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_11_8(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_11_8),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_11_9(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_11_9),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_12_0(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_12_0),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_12_1(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_12_1),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_12_2(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_12_2),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_12_3(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_12_3),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_12_4(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_12_4),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_12_5(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_12_5),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_12_6(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_12_6),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_12_7(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_12_7),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_12_8(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_12_8),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_12_9(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_12_9),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_13_0(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_13_0),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_13_1(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_13_1),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_13_2(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_13_2),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_13_3(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_13_3),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_13_4(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_13_4),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_13_5(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_13_5),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_13_6(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_13_6),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_13_7(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_13_7),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_13_8(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_13_8),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_13_9(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_13_9),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_14_0(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_14_0),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_14_1(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_14_1),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_14_2(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_14_2),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_14_3(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_14_3),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_14_4(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_14_4),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_14_5(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_14_5),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_14_6(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_14_6),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_14_7(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_14_7),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_14_8(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_14_8),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_14_9(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_14_9),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_15_0(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_15_0),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_15_1(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_15_1),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_15_2(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_15_2),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_15_3(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_15_3),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_15_4(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_15_4),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_15_5(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_15_5),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_15_6(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_15_6),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_15_7(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_15_7),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_15_8(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_15_8),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_15_9(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_15_9),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_16_0(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_16_0),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_16_1(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_16_1),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_16_2(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_16_2),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_16_3(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_16_3),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_16_4(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_16_4),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_16_5(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_16_5),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_16_6(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_16_6),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_16_7(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_16_7),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_16_8(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_16_8),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_16_9(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_16_9),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_17_0(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_17_0),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_17_1(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_17_1),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_17_2(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_17_2),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_17_3(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_17_3),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_17_4(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_17_4),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_17_5(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_17_5),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_17_6(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_17_6),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_17_7(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_17_7),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_17_8(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_17_8),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_17_9(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_17_9),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_18_0(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_18_0),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_18_1(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_18_1),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_18_2(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_18_2),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_18_3(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_18_3),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_18_4(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_18_4),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_18_5(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_18_5),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_18_6(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_18_6),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_18_7(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_18_7),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_18_8(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_18_8),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_18_9(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_18_9),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_19_0(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_19_0),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_19_1(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_19_1),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_19_2(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_19_2),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_19_3(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_19_3),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_19_4(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_19_4),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_19_5(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_19_5),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_19_6(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_19_6),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_19_7(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_19_7),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_19_8(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_19_8),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_19_9(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_19_9),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_20_0(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_20_0),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_20_1(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_20_1),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_20_2(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_20_2),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_20_3(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_20_3),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_20_4(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_20_4),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_20_5(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_20_5),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_20_6(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_20_6),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_20_7(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_20_7),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_20_8(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_20_8),
    .io_inConf_bits_confneuralNetsmidAndOutputWeights_20_9(wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_20_9),
    .io_inConf_bits_confneuralNetsbiasVecs_0_0(wellness_io_inConf_bits_confneuralNetsbiasVecs_0_0),
    .io_inConf_bits_confneuralNetsbiasVecs_0_1(wellness_io_inConf_bits_confneuralNetsbiasVecs_0_1),
    .io_inConf_bits_confneuralNetsbiasVecs_0_2(wellness_io_inConf_bits_confneuralNetsbiasVecs_0_2),
    .io_inConf_bits_confneuralNetsbiasVecs_0_3(wellness_io_inConf_bits_confneuralNetsbiasVecs_0_3),
    .io_inConf_bits_confneuralNetsbiasVecs_0_4(wellness_io_inConf_bits_confneuralNetsbiasVecs_0_4),
    .io_inConf_bits_confneuralNetsbiasVecs_0_5(wellness_io_inConf_bits_confneuralNetsbiasVecs_0_5),
    .io_inConf_bits_confneuralNetsbiasVecs_0_6(wellness_io_inConf_bits_confneuralNetsbiasVecs_0_6),
    .io_inConf_bits_confneuralNetsbiasVecs_0_7(wellness_io_inConf_bits_confneuralNetsbiasVecs_0_7),
    .io_inConf_bits_confneuralNetsbiasVecs_0_8(wellness_io_inConf_bits_confneuralNetsbiasVecs_0_8),
    .io_inConf_bits_confneuralNetsbiasVecs_0_9(wellness_io_inConf_bits_confneuralNetsbiasVecs_0_9),
    .io_inConf_bits_confneuralNetsbiasVecs_1_0(wellness_io_inConf_bits_confneuralNetsbiasVecs_1_0),
    .io_inConf_bits_confneuralNetsbiasVecs_1_1(wellness_io_inConf_bits_confneuralNetsbiasVecs_1_1),
    .io_inConf_bits_confneuralNetsbiasVecs_1_2(wellness_io_inConf_bits_confneuralNetsbiasVecs_1_2),
    .io_inConf_bits_confneuralNetsbiasVecs_1_3(wellness_io_inConf_bits_confneuralNetsbiasVecs_1_3),
    .io_inConf_bits_confneuralNetsbiasVecs_1_4(wellness_io_inConf_bits_confneuralNetsbiasVecs_1_4),
    .io_inConf_bits_confneuralNetsbiasVecs_1_5(wellness_io_inConf_bits_confneuralNetsbiasVecs_1_5),
    .io_inConf_bits_confneuralNetsbiasVecs_1_6(wellness_io_inConf_bits_confneuralNetsbiasVecs_1_6),
    .io_inConf_bits_confneuralNetsbiasVecs_1_7(wellness_io_inConf_bits_confneuralNetsbiasVecs_1_7),
    .io_inConf_bits_confneuralNetsbiasVecs_1_8(wellness_io_inConf_bits_confneuralNetsbiasVecs_1_8),
    .io_inConf_bits_confneuralNetsbiasVecs_1_9(wellness_io_inConf_bits_confneuralNetsbiasVecs_1_9),
    .io_inConf_bits_confneuralNetsbiasVecs_2_0(wellness_io_inConf_bits_confneuralNetsbiasVecs_2_0),
    .io_inConf_bits_confneuralNetsbiasVecs_2_1(wellness_io_inConf_bits_confneuralNetsbiasVecs_2_1),
    .io_inConf_bits_confneuralNetsbiasVecs_2_2(wellness_io_inConf_bits_confneuralNetsbiasVecs_2_2),
    .io_inConf_bits_confneuralNetsbiasVecs_2_3(wellness_io_inConf_bits_confneuralNetsbiasVecs_2_3),
    .io_inConf_bits_confneuralNetsbiasVecs_2_4(wellness_io_inConf_bits_confneuralNetsbiasVecs_2_4),
    .io_inConf_bits_confneuralNetsbiasVecs_2_5(wellness_io_inConf_bits_confneuralNetsbiasVecs_2_5),
    .io_inConf_bits_confneuralNetsbiasVecs_2_6(wellness_io_inConf_bits_confneuralNetsbiasVecs_2_6),
    .io_inConf_bits_confneuralNetsbiasVecs_2_7(wellness_io_inConf_bits_confneuralNetsbiasVecs_2_7),
    .io_inConf_bits_confneuralNetsbiasVecs_2_8(wellness_io_inConf_bits_confneuralNetsbiasVecs_2_8),
    .io_inConf_bits_confneuralNetsbiasVecs_2_9(wellness_io_inConf_bits_confneuralNetsbiasVecs_2_9),
    .io_inConf_bits_confneuralNetsoutputBias_0(wellness_io_inConf_bits_confneuralNetsoutputBias_0),
    .io_inConf_bits_confInputMuxSel(wellness_io_inConf_bits_confInputMuxSel),
    .io_out_valid(wellness_io_out_valid),
    .io_out_bits(wellness_io_out_bits),
    .io_rawVotes(wellness_io_rawVotes)
  );
  ConfigurationMemory configurationMemory ( // @[Wellness.scala 398:37]
    .clock(configurationMemory_clock),
    .reset(configurationMemory_reset),
    .io_in_valid(configurationMemory_io_in_valid),
    .io_in_bits_wrdata(configurationMemory_io_in_bits_wrdata),
    .io_in_bits_wraddr(configurationMemory_io_in_bits_wraddr),
    .io_out_bits_confneuralNetsinputWeights_0_0(configurationMemory_io_out_bits_confneuralNetsinputWeights_0_0),
    .io_out_bits_confneuralNetsinputWeights_0_1(configurationMemory_io_out_bits_confneuralNetsinputWeights_0_1),
    .io_out_bits_confneuralNetsinputWeights_0_2(configurationMemory_io_out_bits_confneuralNetsinputWeights_0_2),
    .io_out_bits_confneuralNetsinputWeights_0_3(configurationMemory_io_out_bits_confneuralNetsinputWeights_0_3),
    .io_out_bits_confneuralNetsinputWeights_1_0(configurationMemory_io_out_bits_confneuralNetsinputWeights_1_0),
    .io_out_bits_confneuralNetsinputWeights_1_1(configurationMemory_io_out_bits_confneuralNetsinputWeights_1_1),
    .io_out_bits_confneuralNetsinputWeights_1_2(configurationMemory_io_out_bits_confneuralNetsinputWeights_1_2),
    .io_out_bits_confneuralNetsinputWeights_1_3(configurationMemory_io_out_bits_confneuralNetsinputWeights_1_3),
    .io_out_bits_confneuralNetsinputWeights_2_0(configurationMemory_io_out_bits_confneuralNetsinputWeights_2_0),
    .io_out_bits_confneuralNetsinputWeights_2_1(configurationMemory_io_out_bits_confneuralNetsinputWeights_2_1),
    .io_out_bits_confneuralNetsinputWeights_2_2(configurationMemory_io_out_bits_confneuralNetsinputWeights_2_2),
    .io_out_bits_confneuralNetsinputWeights_2_3(configurationMemory_io_out_bits_confneuralNetsinputWeights_2_3),
    .io_out_bits_confneuralNetsinputWeights_3_0(configurationMemory_io_out_bits_confneuralNetsinputWeights_3_0),
    .io_out_bits_confneuralNetsinputWeights_3_1(configurationMemory_io_out_bits_confneuralNetsinputWeights_3_1),
    .io_out_bits_confneuralNetsinputWeights_3_2(configurationMemory_io_out_bits_confneuralNetsinputWeights_3_2),
    .io_out_bits_confneuralNetsinputWeights_3_3(configurationMemory_io_out_bits_confneuralNetsinputWeights_3_3),
    .io_out_bits_confneuralNetsinputWeights_4_0(configurationMemory_io_out_bits_confneuralNetsinputWeights_4_0),
    .io_out_bits_confneuralNetsinputWeights_4_1(configurationMemory_io_out_bits_confneuralNetsinputWeights_4_1),
    .io_out_bits_confneuralNetsinputWeights_4_2(configurationMemory_io_out_bits_confneuralNetsinputWeights_4_2),
    .io_out_bits_confneuralNetsinputWeights_4_3(configurationMemory_io_out_bits_confneuralNetsinputWeights_4_3),
    .io_out_bits_confneuralNetsinputWeights_5_0(configurationMemory_io_out_bits_confneuralNetsinputWeights_5_0),
    .io_out_bits_confneuralNetsinputWeights_5_1(configurationMemory_io_out_bits_confneuralNetsinputWeights_5_1),
    .io_out_bits_confneuralNetsinputWeights_5_2(configurationMemory_io_out_bits_confneuralNetsinputWeights_5_2),
    .io_out_bits_confneuralNetsinputWeights_5_3(configurationMemory_io_out_bits_confneuralNetsinputWeights_5_3),
    .io_out_bits_confneuralNetsinputWeights_6_0(configurationMemory_io_out_bits_confneuralNetsinputWeights_6_0),
    .io_out_bits_confneuralNetsinputWeights_6_1(configurationMemory_io_out_bits_confneuralNetsinputWeights_6_1),
    .io_out_bits_confneuralNetsinputWeights_6_2(configurationMemory_io_out_bits_confneuralNetsinputWeights_6_2),
    .io_out_bits_confneuralNetsinputWeights_6_3(configurationMemory_io_out_bits_confneuralNetsinputWeights_6_3),
    .io_out_bits_confneuralNetsinputWeights_7_0(configurationMemory_io_out_bits_confneuralNetsinputWeights_7_0),
    .io_out_bits_confneuralNetsinputWeights_7_1(configurationMemory_io_out_bits_confneuralNetsinputWeights_7_1),
    .io_out_bits_confneuralNetsinputWeights_7_2(configurationMemory_io_out_bits_confneuralNetsinputWeights_7_2),
    .io_out_bits_confneuralNetsinputWeights_7_3(configurationMemory_io_out_bits_confneuralNetsinputWeights_7_3),
    .io_out_bits_confneuralNetsinputWeights_8_0(configurationMemory_io_out_bits_confneuralNetsinputWeights_8_0),
    .io_out_bits_confneuralNetsinputWeights_8_1(configurationMemory_io_out_bits_confneuralNetsinputWeights_8_1),
    .io_out_bits_confneuralNetsinputWeights_8_2(configurationMemory_io_out_bits_confneuralNetsinputWeights_8_2),
    .io_out_bits_confneuralNetsinputWeights_8_3(configurationMemory_io_out_bits_confneuralNetsinputWeights_8_3),
    .io_out_bits_confneuralNetsinputWeights_9_0(configurationMemory_io_out_bits_confneuralNetsinputWeights_9_0),
    .io_out_bits_confneuralNetsinputWeights_9_1(configurationMemory_io_out_bits_confneuralNetsinputWeights_9_1),
    .io_out_bits_confneuralNetsinputWeights_9_2(configurationMemory_io_out_bits_confneuralNetsinputWeights_9_2),
    .io_out_bits_confneuralNetsinputWeights_9_3(configurationMemory_io_out_bits_confneuralNetsinputWeights_9_3),
    .io_out_bits_confneuralNetsmidAndOutputWeights_0_0(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_0_0),
    .io_out_bits_confneuralNetsmidAndOutputWeights_0_1(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_0_1),
    .io_out_bits_confneuralNetsmidAndOutputWeights_0_2(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_0_2),
    .io_out_bits_confneuralNetsmidAndOutputWeights_0_3(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_0_3),
    .io_out_bits_confneuralNetsmidAndOutputWeights_0_4(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_0_4),
    .io_out_bits_confneuralNetsmidAndOutputWeights_0_5(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_0_5),
    .io_out_bits_confneuralNetsmidAndOutputWeights_0_6(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_0_6),
    .io_out_bits_confneuralNetsmidAndOutputWeights_0_7(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_0_7),
    .io_out_bits_confneuralNetsmidAndOutputWeights_0_8(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_0_8),
    .io_out_bits_confneuralNetsmidAndOutputWeights_0_9(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_0_9),
    .io_out_bits_confneuralNetsmidAndOutputWeights_1_0(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_1_0),
    .io_out_bits_confneuralNetsmidAndOutputWeights_1_1(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_1_1),
    .io_out_bits_confneuralNetsmidAndOutputWeights_1_2(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_1_2),
    .io_out_bits_confneuralNetsmidAndOutputWeights_1_3(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_1_3),
    .io_out_bits_confneuralNetsmidAndOutputWeights_1_4(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_1_4),
    .io_out_bits_confneuralNetsmidAndOutputWeights_1_5(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_1_5),
    .io_out_bits_confneuralNetsmidAndOutputWeights_1_6(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_1_6),
    .io_out_bits_confneuralNetsmidAndOutputWeights_1_7(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_1_7),
    .io_out_bits_confneuralNetsmidAndOutputWeights_1_8(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_1_8),
    .io_out_bits_confneuralNetsmidAndOutputWeights_1_9(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_1_9),
    .io_out_bits_confneuralNetsmidAndOutputWeights_2_0(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_2_0),
    .io_out_bits_confneuralNetsmidAndOutputWeights_2_1(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_2_1),
    .io_out_bits_confneuralNetsmidAndOutputWeights_2_2(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_2_2),
    .io_out_bits_confneuralNetsmidAndOutputWeights_2_3(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_2_3),
    .io_out_bits_confneuralNetsmidAndOutputWeights_2_4(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_2_4),
    .io_out_bits_confneuralNetsmidAndOutputWeights_2_5(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_2_5),
    .io_out_bits_confneuralNetsmidAndOutputWeights_2_6(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_2_6),
    .io_out_bits_confneuralNetsmidAndOutputWeights_2_7(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_2_7),
    .io_out_bits_confneuralNetsmidAndOutputWeights_2_8(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_2_8),
    .io_out_bits_confneuralNetsmidAndOutputWeights_2_9(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_2_9),
    .io_out_bits_confneuralNetsmidAndOutputWeights_3_0(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_3_0),
    .io_out_bits_confneuralNetsmidAndOutputWeights_3_1(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_3_1),
    .io_out_bits_confneuralNetsmidAndOutputWeights_3_2(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_3_2),
    .io_out_bits_confneuralNetsmidAndOutputWeights_3_3(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_3_3),
    .io_out_bits_confneuralNetsmidAndOutputWeights_3_4(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_3_4),
    .io_out_bits_confneuralNetsmidAndOutputWeights_3_5(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_3_5),
    .io_out_bits_confneuralNetsmidAndOutputWeights_3_6(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_3_6),
    .io_out_bits_confneuralNetsmidAndOutputWeights_3_7(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_3_7),
    .io_out_bits_confneuralNetsmidAndOutputWeights_3_8(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_3_8),
    .io_out_bits_confneuralNetsmidAndOutputWeights_3_9(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_3_9),
    .io_out_bits_confneuralNetsmidAndOutputWeights_4_0(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_4_0),
    .io_out_bits_confneuralNetsmidAndOutputWeights_4_1(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_4_1),
    .io_out_bits_confneuralNetsmidAndOutputWeights_4_2(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_4_2),
    .io_out_bits_confneuralNetsmidAndOutputWeights_4_3(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_4_3),
    .io_out_bits_confneuralNetsmidAndOutputWeights_4_4(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_4_4),
    .io_out_bits_confneuralNetsmidAndOutputWeights_4_5(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_4_5),
    .io_out_bits_confneuralNetsmidAndOutputWeights_4_6(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_4_6),
    .io_out_bits_confneuralNetsmidAndOutputWeights_4_7(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_4_7),
    .io_out_bits_confneuralNetsmidAndOutputWeights_4_8(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_4_8),
    .io_out_bits_confneuralNetsmidAndOutputWeights_4_9(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_4_9),
    .io_out_bits_confneuralNetsmidAndOutputWeights_5_0(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_5_0),
    .io_out_bits_confneuralNetsmidAndOutputWeights_5_1(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_5_1),
    .io_out_bits_confneuralNetsmidAndOutputWeights_5_2(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_5_2),
    .io_out_bits_confneuralNetsmidAndOutputWeights_5_3(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_5_3),
    .io_out_bits_confneuralNetsmidAndOutputWeights_5_4(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_5_4),
    .io_out_bits_confneuralNetsmidAndOutputWeights_5_5(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_5_5),
    .io_out_bits_confneuralNetsmidAndOutputWeights_5_6(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_5_6),
    .io_out_bits_confneuralNetsmidAndOutputWeights_5_7(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_5_7),
    .io_out_bits_confneuralNetsmidAndOutputWeights_5_8(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_5_8),
    .io_out_bits_confneuralNetsmidAndOutputWeights_5_9(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_5_9),
    .io_out_bits_confneuralNetsmidAndOutputWeights_6_0(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_6_0),
    .io_out_bits_confneuralNetsmidAndOutputWeights_6_1(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_6_1),
    .io_out_bits_confneuralNetsmidAndOutputWeights_6_2(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_6_2),
    .io_out_bits_confneuralNetsmidAndOutputWeights_6_3(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_6_3),
    .io_out_bits_confneuralNetsmidAndOutputWeights_6_4(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_6_4),
    .io_out_bits_confneuralNetsmidAndOutputWeights_6_5(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_6_5),
    .io_out_bits_confneuralNetsmidAndOutputWeights_6_6(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_6_6),
    .io_out_bits_confneuralNetsmidAndOutputWeights_6_7(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_6_7),
    .io_out_bits_confneuralNetsmidAndOutputWeights_6_8(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_6_8),
    .io_out_bits_confneuralNetsmidAndOutputWeights_6_9(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_6_9),
    .io_out_bits_confneuralNetsmidAndOutputWeights_7_0(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_7_0),
    .io_out_bits_confneuralNetsmidAndOutputWeights_7_1(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_7_1),
    .io_out_bits_confneuralNetsmidAndOutputWeights_7_2(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_7_2),
    .io_out_bits_confneuralNetsmidAndOutputWeights_7_3(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_7_3),
    .io_out_bits_confneuralNetsmidAndOutputWeights_7_4(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_7_4),
    .io_out_bits_confneuralNetsmidAndOutputWeights_7_5(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_7_5),
    .io_out_bits_confneuralNetsmidAndOutputWeights_7_6(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_7_6),
    .io_out_bits_confneuralNetsmidAndOutputWeights_7_7(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_7_7),
    .io_out_bits_confneuralNetsmidAndOutputWeights_7_8(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_7_8),
    .io_out_bits_confneuralNetsmidAndOutputWeights_7_9(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_7_9),
    .io_out_bits_confneuralNetsmidAndOutputWeights_8_0(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_8_0),
    .io_out_bits_confneuralNetsmidAndOutputWeights_8_1(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_8_1),
    .io_out_bits_confneuralNetsmidAndOutputWeights_8_2(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_8_2),
    .io_out_bits_confneuralNetsmidAndOutputWeights_8_3(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_8_3),
    .io_out_bits_confneuralNetsmidAndOutputWeights_8_4(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_8_4),
    .io_out_bits_confneuralNetsmidAndOutputWeights_8_5(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_8_5),
    .io_out_bits_confneuralNetsmidAndOutputWeights_8_6(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_8_6),
    .io_out_bits_confneuralNetsmidAndOutputWeights_8_7(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_8_7),
    .io_out_bits_confneuralNetsmidAndOutputWeights_8_8(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_8_8),
    .io_out_bits_confneuralNetsmidAndOutputWeights_8_9(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_8_9),
    .io_out_bits_confneuralNetsmidAndOutputWeights_9_0(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_9_0),
    .io_out_bits_confneuralNetsmidAndOutputWeights_9_1(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_9_1),
    .io_out_bits_confneuralNetsmidAndOutputWeights_9_2(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_9_2),
    .io_out_bits_confneuralNetsmidAndOutputWeights_9_3(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_9_3),
    .io_out_bits_confneuralNetsmidAndOutputWeights_9_4(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_9_4),
    .io_out_bits_confneuralNetsmidAndOutputWeights_9_5(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_9_5),
    .io_out_bits_confneuralNetsmidAndOutputWeights_9_6(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_9_6),
    .io_out_bits_confneuralNetsmidAndOutputWeights_9_7(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_9_7),
    .io_out_bits_confneuralNetsmidAndOutputWeights_9_8(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_9_8),
    .io_out_bits_confneuralNetsmidAndOutputWeights_9_9(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_9_9),
    .io_out_bits_confneuralNetsmidAndOutputWeights_10_0(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_10_0),
    .io_out_bits_confneuralNetsmidAndOutputWeights_10_1(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_10_1),
    .io_out_bits_confneuralNetsmidAndOutputWeights_10_2(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_10_2),
    .io_out_bits_confneuralNetsmidAndOutputWeights_10_3(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_10_3),
    .io_out_bits_confneuralNetsmidAndOutputWeights_10_4(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_10_4),
    .io_out_bits_confneuralNetsmidAndOutputWeights_10_5(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_10_5),
    .io_out_bits_confneuralNetsmidAndOutputWeights_10_6(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_10_6),
    .io_out_bits_confneuralNetsmidAndOutputWeights_10_7(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_10_7),
    .io_out_bits_confneuralNetsmidAndOutputWeights_10_8(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_10_8),
    .io_out_bits_confneuralNetsmidAndOutputWeights_10_9(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_10_9),
    .io_out_bits_confneuralNetsmidAndOutputWeights_11_0(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_11_0),
    .io_out_bits_confneuralNetsmidAndOutputWeights_11_1(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_11_1),
    .io_out_bits_confneuralNetsmidAndOutputWeights_11_2(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_11_2),
    .io_out_bits_confneuralNetsmidAndOutputWeights_11_3(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_11_3),
    .io_out_bits_confneuralNetsmidAndOutputWeights_11_4(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_11_4),
    .io_out_bits_confneuralNetsmidAndOutputWeights_11_5(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_11_5),
    .io_out_bits_confneuralNetsmidAndOutputWeights_11_6(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_11_6),
    .io_out_bits_confneuralNetsmidAndOutputWeights_11_7(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_11_7),
    .io_out_bits_confneuralNetsmidAndOutputWeights_11_8(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_11_8),
    .io_out_bits_confneuralNetsmidAndOutputWeights_11_9(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_11_9),
    .io_out_bits_confneuralNetsmidAndOutputWeights_12_0(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_12_0),
    .io_out_bits_confneuralNetsmidAndOutputWeights_12_1(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_12_1),
    .io_out_bits_confneuralNetsmidAndOutputWeights_12_2(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_12_2),
    .io_out_bits_confneuralNetsmidAndOutputWeights_12_3(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_12_3),
    .io_out_bits_confneuralNetsmidAndOutputWeights_12_4(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_12_4),
    .io_out_bits_confneuralNetsmidAndOutputWeights_12_5(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_12_5),
    .io_out_bits_confneuralNetsmidAndOutputWeights_12_6(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_12_6),
    .io_out_bits_confneuralNetsmidAndOutputWeights_12_7(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_12_7),
    .io_out_bits_confneuralNetsmidAndOutputWeights_12_8(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_12_8),
    .io_out_bits_confneuralNetsmidAndOutputWeights_12_9(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_12_9),
    .io_out_bits_confneuralNetsmidAndOutputWeights_13_0(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_13_0),
    .io_out_bits_confneuralNetsmidAndOutputWeights_13_1(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_13_1),
    .io_out_bits_confneuralNetsmidAndOutputWeights_13_2(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_13_2),
    .io_out_bits_confneuralNetsmidAndOutputWeights_13_3(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_13_3),
    .io_out_bits_confneuralNetsmidAndOutputWeights_13_4(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_13_4),
    .io_out_bits_confneuralNetsmidAndOutputWeights_13_5(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_13_5),
    .io_out_bits_confneuralNetsmidAndOutputWeights_13_6(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_13_6),
    .io_out_bits_confneuralNetsmidAndOutputWeights_13_7(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_13_7),
    .io_out_bits_confneuralNetsmidAndOutputWeights_13_8(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_13_8),
    .io_out_bits_confneuralNetsmidAndOutputWeights_13_9(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_13_9),
    .io_out_bits_confneuralNetsmidAndOutputWeights_14_0(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_14_0),
    .io_out_bits_confneuralNetsmidAndOutputWeights_14_1(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_14_1),
    .io_out_bits_confneuralNetsmidAndOutputWeights_14_2(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_14_2),
    .io_out_bits_confneuralNetsmidAndOutputWeights_14_3(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_14_3),
    .io_out_bits_confneuralNetsmidAndOutputWeights_14_4(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_14_4),
    .io_out_bits_confneuralNetsmidAndOutputWeights_14_5(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_14_5),
    .io_out_bits_confneuralNetsmidAndOutputWeights_14_6(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_14_6),
    .io_out_bits_confneuralNetsmidAndOutputWeights_14_7(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_14_7),
    .io_out_bits_confneuralNetsmidAndOutputWeights_14_8(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_14_8),
    .io_out_bits_confneuralNetsmidAndOutputWeights_14_9(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_14_9),
    .io_out_bits_confneuralNetsmidAndOutputWeights_15_0(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_15_0),
    .io_out_bits_confneuralNetsmidAndOutputWeights_15_1(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_15_1),
    .io_out_bits_confneuralNetsmidAndOutputWeights_15_2(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_15_2),
    .io_out_bits_confneuralNetsmidAndOutputWeights_15_3(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_15_3),
    .io_out_bits_confneuralNetsmidAndOutputWeights_15_4(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_15_4),
    .io_out_bits_confneuralNetsmidAndOutputWeights_15_5(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_15_5),
    .io_out_bits_confneuralNetsmidAndOutputWeights_15_6(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_15_6),
    .io_out_bits_confneuralNetsmidAndOutputWeights_15_7(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_15_7),
    .io_out_bits_confneuralNetsmidAndOutputWeights_15_8(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_15_8),
    .io_out_bits_confneuralNetsmidAndOutputWeights_15_9(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_15_9),
    .io_out_bits_confneuralNetsmidAndOutputWeights_16_0(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_16_0),
    .io_out_bits_confneuralNetsmidAndOutputWeights_16_1(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_16_1),
    .io_out_bits_confneuralNetsmidAndOutputWeights_16_2(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_16_2),
    .io_out_bits_confneuralNetsmidAndOutputWeights_16_3(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_16_3),
    .io_out_bits_confneuralNetsmidAndOutputWeights_16_4(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_16_4),
    .io_out_bits_confneuralNetsmidAndOutputWeights_16_5(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_16_5),
    .io_out_bits_confneuralNetsmidAndOutputWeights_16_6(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_16_6),
    .io_out_bits_confneuralNetsmidAndOutputWeights_16_7(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_16_7),
    .io_out_bits_confneuralNetsmidAndOutputWeights_16_8(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_16_8),
    .io_out_bits_confneuralNetsmidAndOutputWeights_16_9(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_16_9),
    .io_out_bits_confneuralNetsmidAndOutputWeights_17_0(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_17_0),
    .io_out_bits_confneuralNetsmidAndOutputWeights_17_1(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_17_1),
    .io_out_bits_confneuralNetsmidAndOutputWeights_17_2(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_17_2),
    .io_out_bits_confneuralNetsmidAndOutputWeights_17_3(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_17_3),
    .io_out_bits_confneuralNetsmidAndOutputWeights_17_4(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_17_4),
    .io_out_bits_confneuralNetsmidAndOutputWeights_17_5(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_17_5),
    .io_out_bits_confneuralNetsmidAndOutputWeights_17_6(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_17_6),
    .io_out_bits_confneuralNetsmidAndOutputWeights_17_7(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_17_7),
    .io_out_bits_confneuralNetsmidAndOutputWeights_17_8(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_17_8),
    .io_out_bits_confneuralNetsmidAndOutputWeights_17_9(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_17_9),
    .io_out_bits_confneuralNetsmidAndOutputWeights_18_0(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_18_0),
    .io_out_bits_confneuralNetsmidAndOutputWeights_18_1(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_18_1),
    .io_out_bits_confneuralNetsmidAndOutputWeights_18_2(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_18_2),
    .io_out_bits_confneuralNetsmidAndOutputWeights_18_3(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_18_3),
    .io_out_bits_confneuralNetsmidAndOutputWeights_18_4(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_18_4),
    .io_out_bits_confneuralNetsmidAndOutputWeights_18_5(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_18_5),
    .io_out_bits_confneuralNetsmidAndOutputWeights_18_6(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_18_6),
    .io_out_bits_confneuralNetsmidAndOutputWeights_18_7(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_18_7),
    .io_out_bits_confneuralNetsmidAndOutputWeights_18_8(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_18_8),
    .io_out_bits_confneuralNetsmidAndOutputWeights_18_9(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_18_9),
    .io_out_bits_confneuralNetsmidAndOutputWeights_19_0(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_19_0),
    .io_out_bits_confneuralNetsmidAndOutputWeights_19_1(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_19_1),
    .io_out_bits_confneuralNetsmidAndOutputWeights_19_2(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_19_2),
    .io_out_bits_confneuralNetsmidAndOutputWeights_19_3(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_19_3),
    .io_out_bits_confneuralNetsmidAndOutputWeights_19_4(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_19_4),
    .io_out_bits_confneuralNetsmidAndOutputWeights_19_5(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_19_5),
    .io_out_bits_confneuralNetsmidAndOutputWeights_19_6(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_19_6),
    .io_out_bits_confneuralNetsmidAndOutputWeights_19_7(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_19_7),
    .io_out_bits_confneuralNetsmidAndOutputWeights_19_8(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_19_8),
    .io_out_bits_confneuralNetsmidAndOutputWeights_19_9(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_19_9),
    .io_out_bits_confneuralNetsmidAndOutputWeights_20_0(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_20_0),
    .io_out_bits_confneuralNetsmidAndOutputWeights_20_1(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_20_1),
    .io_out_bits_confneuralNetsmidAndOutputWeights_20_2(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_20_2),
    .io_out_bits_confneuralNetsmidAndOutputWeights_20_3(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_20_3),
    .io_out_bits_confneuralNetsmidAndOutputWeights_20_4(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_20_4),
    .io_out_bits_confneuralNetsmidAndOutputWeights_20_5(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_20_5),
    .io_out_bits_confneuralNetsmidAndOutputWeights_20_6(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_20_6),
    .io_out_bits_confneuralNetsmidAndOutputWeights_20_7(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_20_7),
    .io_out_bits_confneuralNetsmidAndOutputWeights_20_8(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_20_8),
    .io_out_bits_confneuralNetsmidAndOutputWeights_20_9(configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_20_9),
    .io_out_bits_confneuralNetsbiasVecs_0_0(configurationMemory_io_out_bits_confneuralNetsbiasVecs_0_0),
    .io_out_bits_confneuralNetsbiasVecs_0_1(configurationMemory_io_out_bits_confneuralNetsbiasVecs_0_1),
    .io_out_bits_confneuralNetsbiasVecs_0_2(configurationMemory_io_out_bits_confneuralNetsbiasVecs_0_2),
    .io_out_bits_confneuralNetsbiasVecs_0_3(configurationMemory_io_out_bits_confneuralNetsbiasVecs_0_3),
    .io_out_bits_confneuralNetsbiasVecs_0_4(configurationMemory_io_out_bits_confneuralNetsbiasVecs_0_4),
    .io_out_bits_confneuralNetsbiasVecs_0_5(configurationMemory_io_out_bits_confneuralNetsbiasVecs_0_5),
    .io_out_bits_confneuralNetsbiasVecs_0_6(configurationMemory_io_out_bits_confneuralNetsbiasVecs_0_6),
    .io_out_bits_confneuralNetsbiasVecs_0_7(configurationMemory_io_out_bits_confneuralNetsbiasVecs_0_7),
    .io_out_bits_confneuralNetsbiasVecs_0_8(configurationMemory_io_out_bits_confneuralNetsbiasVecs_0_8),
    .io_out_bits_confneuralNetsbiasVecs_0_9(configurationMemory_io_out_bits_confneuralNetsbiasVecs_0_9),
    .io_out_bits_confneuralNetsbiasVecs_1_0(configurationMemory_io_out_bits_confneuralNetsbiasVecs_1_0),
    .io_out_bits_confneuralNetsbiasVecs_1_1(configurationMemory_io_out_bits_confneuralNetsbiasVecs_1_1),
    .io_out_bits_confneuralNetsbiasVecs_1_2(configurationMemory_io_out_bits_confneuralNetsbiasVecs_1_2),
    .io_out_bits_confneuralNetsbiasVecs_1_3(configurationMemory_io_out_bits_confneuralNetsbiasVecs_1_3),
    .io_out_bits_confneuralNetsbiasVecs_1_4(configurationMemory_io_out_bits_confneuralNetsbiasVecs_1_4),
    .io_out_bits_confneuralNetsbiasVecs_1_5(configurationMemory_io_out_bits_confneuralNetsbiasVecs_1_5),
    .io_out_bits_confneuralNetsbiasVecs_1_6(configurationMemory_io_out_bits_confneuralNetsbiasVecs_1_6),
    .io_out_bits_confneuralNetsbiasVecs_1_7(configurationMemory_io_out_bits_confneuralNetsbiasVecs_1_7),
    .io_out_bits_confneuralNetsbiasVecs_1_8(configurationMemory_io_out_bits_confneuralNetsbiasVecs_1_8),
    .io_out_bits_confneuralNetsbiasVecs_1_9(configurationMemory_io_out_bits_confneuralNetsbiasVecs_1_9),
    .io_out_bits_confneuralNetsbiasVecs_2_0(configurationMemory_io_out_bits_confneuralNetsbiasVecs_2_0),
    .io_out_bits_confneuralNetsbiasVecs_2_1(configurationMemory_io_out_bits_confneuralNetsbiasVecs_2_1),
    .io_out_bits_confneuralNetsbiasVecs_2_2(configurationMemory_io_out_bits_confneuralNetsbiasVecs_2_2),
    .io_out_bits_confneuralNetsbiasVecs_2_3(configurationMemory_io_out_bits_confneuralNetsbiasVecs_2_3),
    .io_out_bits_confneuralNetsbiasVecs_2_4(configurationMemory_io_out_bits_confneuralNetsbiasVecs_2_4),
    .io_out_bits_confneuralNetsbiasVecs_2_5(configurationMemory_io_out_bits_confneuralNetsbiasVecs_2_5),
    .io_out_bits_confneuralNetsbiasVecs_2_6(configurationMemory_io_out_bits_confneuralNetsbiasVecs_2_6),
    .io_out_bits_confneuralNetsbiasVecs_2_7(configurationMemory_io_out_bits_confneuralNetsbiasVecs_2_7),
    .io_out_bits_confneuralNetsbiasVecs_2_8(configurationMemory_io_out_bits_confneuralNetsbiasVecs_2_8),
    .io_out_bits_confneuralNetsbiasVecs_2_9(configurationMemory_io_out_bits_confneuralNetsbiasVecs_2_9),
    .io_out_bits_confneuralNetsoutputBias_0(configurationMemory_io_out_bits_confneuralNetsoutputBias_0),
    .io_out_bits_confInputMuxSel(configurationMemory_io_out_bits_confInputMuxSel)
  );
  assign in_1_bits_data = converter_1_auto_out_bits_data; // @[Nodes.scala 333:76 LazyModule.scala 167:31]
  assign _T_4 = $signed(in_1_bits_data); // @[Wellness.scala 408:49]
  assign _T_5 = $unsigned(wellness_io_rawVotes); // @[Wellness.scala 411:83]
  assign _T_6 = {wellness_io_out_bits,_T_5}; // @[Cat.scala 30:58]
  assign inConf_bits_data = converter_2_auto_out_bits_data; // @[Nodes.scala 333:76 LazyModule.scala 167:31]
  assign _T_7 = inConf_bits_data[31:0]; // @[Wellness.scala 418:62]
  assign _GEN_0 = _T_4[31:0]; // @[Wellness.scala 408:49 Wellness.scala 408:49]
  assign in_ready = converter_1_auto_in_ready; // @[BundleBridge.scala 39:12]
  assign out_valid = converter_auto_out_valid; // @[BundleBridge.scala 27:8]
  assign out_bits_data = converter_auto_out_bits_data; // @[BundleBridge.scala 27:8]
  assign out_bits_last = converter_auto_out_bits_last; // @[BundleBridge.scala 27:8]
  assign in2_ready = converter_2_auto_in_ready; // @[BundleBridge.scala 39:12]
  assign converter_auto_in_valid = wellness_io_out_valid; // @[LazyModule.scala 167:57]
  assign converter_auto_in_bits_data = {{31'd0}, _T_6}; // @[LazyModule.scala 167:57]
  assign converter_auto_in_bits_last = 1'h0; // @[LazyModule.scala 167:57]
  assign converter_auto_out_ready = out_ready; // @[LazyModule.scala 167:31]
  assign converter_1_auto_in_valid = in_valid; // @[LazyModule.scala 167:57]
  assign converter_1_auto_in_bits_data = in_bits_data; // @[LazyModule.scala 167:57]
  assign converter_1_auto_in_bits_last = in_bits_last; // @[LazyModule.scala 167:57]
  assign converter_1_auto_out_ready = 1'h1; // @[LazyModule.scala 167:31]
  assign converter_2_auto_in_valid = in2_valid; // @[LazyModule.scala 167:57]
  assign converter_2_auto_in_bits_data = in2_bits_data; // @[LazyModule.scala 167:57]
  assign converter_2_auto_in_bits_last = in2_bits_last; // @[LazyModule.scala 167:57]
  assign converter_2_auto_out_ready = 1'h1; // @[LazyModule.scala 167:31]
  assign wellness_clock = clock;
  assign wellness_reset = reset;
  assign wellness_io_streamIn_valid = streamIn_valid; // @[Wellness.scala 402:32]
  assign wellness_io_streamIn_bits = streamIn_bits; // @[Wellness.scala 401:31]
  assign wellness_io_in_valid = converter_1_auto_out_valid; // @[Wellness.scala 407:26]
  assign wellness_io_in_bits = $signed(_GEN_0); // @[Wellness.scala 408:25]
  assign wellness_io_inConf_bits_confneuralNetsinputWeights_0_0 = configurationMemory_io_out_bits_confneuralNetsinputWeights_0_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsinputWeights_0_1 = configurationMemory_io_out_bits_confneuralNetsinputWeights_0_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsinputWeights_0_2 = configurationMemory_io_out_bits_confneuralNetsinputWeights_0_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsinputWeights_0_3 = configurationMemory_io_out_bits_confneuralNetsinputWeights_0_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsinputWeights_1_0 = configurationMemory_io_out_bits_confneuralNetsinputWeights_1_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsinputWeights_1_1 = configurationMemory_io_out_bits_confneuralNetsinputWeights_1_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsinputWeights_1_2 = configurationMemory_io_out_bits_confneuralNetsinputWeights_1_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsinputWeights_1_3 = configurationMemory_io_out_bits_confneuralNetsinputWeights_1_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsinputWeights_2_0 = configurationMemory_io_out_bits_confneuralNetsinputWeights_2_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsinputWeights_2_1 = configurationMemory_io_out_bits_confneuralNetsinputWeights_2_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsinputWeights_2_2 = configurationMemory_io_out_bits_confneuralNetsinputWeights_2_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsinputWeights_2_3 = configurationMemory_io_out_bits_confneuralNetsinputWeights_2_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsinputWeights_3_0 = configurationMemory_io_out_bits_confneuralNetsinputWeights_3_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsinputWeights_3_1 = configurationMemory_io_out_bits_confneuralNetsinputWeights_3_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsinputWeights_3_2 = configurationMemory_io_out_bits_confneuralNetsinputWeights_3_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsinputWeights_3_3 = configurationMemory_io_out_bits_confneuralNetsinputWeights_3_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsinputWeights_4_0 = configurationMemory_io_out_bits_confneuralNetsinputWeights_4_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsinputWeights_4_1 = configurationMemory_io_out_bits_confneuralNetsinputWeights_4_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsinputWeights_4_2 = configurationMemory_io_out_bits_confneuralNetsinputWeights_4_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsinputWeights_4_3 = configurationMemory_io_out_bits_confneuralNetsinputWeights_4_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsinputWeights_5_0 = configurationMemory_io_out_bits_confneuralNetsinputWeights_5_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsinputWeights_5_1 = configurationMemory_io_out_bits_confneuralNetsinputWeights_5_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsinputWeights_5_2 = configurationMemory_io_out_bits_confneuralNetsinputWeights_5_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsinputWeights_5_3 = configurationMemory_io_out_bits_confneuralNetsinputWeights_5_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsinputWeights_6_0 = configurationMemory_io_out_bits_confneuralNetsinputWeights_6_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsinputWeights_6_1 = configurationMemory_io_out_bits_confneuralNetsinputWeights_6_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsinputWeights_6_2 = configurationMemory_io_out_bits_confneuralNetsinputWeights_6_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsinputWeights_6_3 = configurationMemory_io_out_bits_confneuralNetsinputWeights_6_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsinputWeights_7_0 = configurationMemory_io_out_bits_confneuralNetsinputWeights_7_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsinputWeights_7_1 = configurationMemory_io_out_bits_confneuralNetsinputWeights_7_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsinputWeights_7_2 = configurationMemory_io_out_bits_confneuralNetsinputWeights_7_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsinputWeights_7_3 = configurationMemory_io_out_bits_confneuralNetsinputWeights_7_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsinputWeights_8_0 = configurationMemory_io_out_bits_confneuralNetsinputWeights_8_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsinputWeights_8_1 = configurationMemory_io_out_bits_confneuralNetsinputWeights_8_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsinputWeights_8_2 = configurationMemory_io_out_bits_confneuralNetsinputWeights_8_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsinputWeights_8_3 = configurationMemory_io_out_bits_confneuralNetsinputWeights_8_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsinputWeights_9_0 = configurationMemory_io_out_bits_confneuralNetsinputWeights_9_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsinputWeights_9_1 = configurationMemory_io_out_bits_confneuralNetsinputWeights_9_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsinputWeights_9_2 = configurationMemory_io_out_bits_confneuralNetsinputWeights_9_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsinputWeights_9_3 = configurationMemory_io_out_bits_confneuralNetsinputWeights_9_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_0_0 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_0_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_0_1 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_0_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_0_2 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_0_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_0_3 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_0_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_0_4 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_0_4; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_0_5 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_0_5; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_0_6 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_0_6; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_0_7 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_0_7; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_0_8 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_0_8; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_0_9 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_0_9; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_1_0 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_1_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_1_1 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_1_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_1_2 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_1_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_1_3 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_1_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_1_4 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_1_4; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_1_5 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_1_5; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_1_6 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_1_6; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_1_7 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_1_7; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_1_8 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_1_8; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_1_9 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_1_9; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_2_0 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_2_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_2_1 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_2_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_2_2 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_2_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_2_3 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_2_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_2_4 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_2_4; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_2_5 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_2_5; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_2_6 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_2_6; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_2_7 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_2_7; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_2_8 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_2_8; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_2_9 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_2_9; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_3_0 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_3_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_3_1 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_3_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_3_2 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_3_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_3_3 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_3_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_3_4 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_3_4; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_3_5 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_3_5; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_3_6 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_3_6; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_3_7 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_3_7; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_3_8 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_3_8; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_3_9 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_3_9; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_4_0 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_4_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_4_1 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_4_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_4_2 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_4_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_4_3 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_4_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_4_4 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_4_4; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_4_5 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_4_5; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_4_6 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_4_6; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_4_7 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_4_7; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_4_8 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_4_8; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_4_9 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_4_9; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_5_0 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_5_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_5_1 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_5_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_5_2 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_5_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_5_3 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_5_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_5_4 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_5_4; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_5_5 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_5_5; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_5_6 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_5_6; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_5_7 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_5_7; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_5_8 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_5_8; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_5_9 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_5_9; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_6_0 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_6_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_6_1 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_6_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_6_2 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_6_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_6_3 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_6_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_6_4 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_6_4; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_6_5 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_6_5; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_6_6 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_6_6; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_6_7 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_6_7; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_6_8 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_6_8; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_6_9 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_6_9; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_7_0 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_7_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_7_1 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_7_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_7_2 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_7_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_7_3 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_7_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_7_4 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_7_4; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_7_5 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_7_5; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_7_6 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_7_6; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_7_7 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_7_7; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_7_8 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_7_8; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_7_9 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_7_9; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_8_0 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_8_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_8_1 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_8_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_8_2 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_8_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_8_3 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_8_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_8_4 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_8_4; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_8_5 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_8_5; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_8_6 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_8_6; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_8_7 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_8_7; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_8_8 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_8_8; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_8_9 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_8_9; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_9_0 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_9_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_9_1 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_9_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_9_2 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_9_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_9_3 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_9_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_9_4 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_9_4; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_9_5 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_9_5; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_9_6 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_9_6; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_9_7 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_9_7; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_9_8 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_9_8; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_9_9 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_9_9; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_10_0 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_10_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_10_1 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_10_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_10_2 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_10_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_10_3 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_10_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_10_4 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_10_4; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_10_5 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_10_5; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_10_6 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_10_6; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_10_7 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_10_7; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_10_8 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_10_8; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_10_9 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_10_9; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_11_0 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_11_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_11_1 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_11_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_11_2 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_11_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_11_3 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_11_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_11_4 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_11_4; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_11_5 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_11_5; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_11_6 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_11_6; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_11_7 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_11_7; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_11_8 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_11_8; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_11_9 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_11_9; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_12_0 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_12_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_12_1 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_12_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_12_2 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_12_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_12_3 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_12_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_12_4 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_12_4; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_12_5 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_12_5; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_12_6 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_12_6; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_12_7 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_12_7; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_12_8 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_12_8; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_12_9 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_12_9; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_13_0 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_13_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_13_1 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_13_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_13_2 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_13_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_13_3 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_13_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_13_4 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_13_4; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_13_5 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_13_5; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_13_6 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_13_6; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_13_7 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_13_7; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_13_8 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_13_8; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_13_9 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_13_9; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_14_0 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_14_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_14_1 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_14_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_14_2 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_14_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_14_3 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_14_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_14_4 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_14_4; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_14_5 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_14_5; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_14_6 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_14_6; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_14_7 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_14_7; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_14_8 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_14_8; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_14_9 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_14_9; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_15_0 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_15_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_15_1 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_15_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_15_2 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_15_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_15_3 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_15_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_15_4 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_15_4; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_15_5 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_15_5; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_15_6 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_15_6; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_15_7 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_15_7; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_15_8 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_15_8; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_15_9 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_15_9; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_16_0 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_16_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_16_1 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_16_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_16_2 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_16_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_16_3 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_16_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_16_4 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_16_4; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_16_5 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_16_5; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_16_6 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_16_6; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_16_7 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_16_7; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_16_8 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_16_8; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_16_9 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_16_9; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_17_0 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_17_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_17_1 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_17_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_17_2 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_17_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_17_3 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_17_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_17_4 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_17_4; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_17_5 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_17_5; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_17_6 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_17_6; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_17_7 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_17_7; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_17_8 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_17_8; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_17_9 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_17_9; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_18_0 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_18_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_18_1 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_18_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_18_2 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_18_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_18_3 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_18_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_18_4 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_18_4; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_18_5 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_18_5; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_18_6 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_18_6; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_18_7 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_18_7; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_18_8 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_18_8; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_18_9 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_18_9; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_19_0 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_19_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_19_1 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_19_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_19_2 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_19_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_19_3 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_19_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_19_4 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_19_4; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_19_5 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_19_5; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_19_6 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_19_6; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_19_7 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_19_7; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_19_8 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_19_8; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_19_9 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_19_9; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_20_0 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_20_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_20_1 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_20_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_20_2 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_20_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_20_3 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_20_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_20_4 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_20_4; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_20_5 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_20_5; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_20_6 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_20_6; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_20_7 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_20_7; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_20_8 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_20_8; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsmidAndOutputWeights_20_9 = configurationMemory_io_out_bits_confneuralNetsmidAndOutputWeights_20_9; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVecs_0_0 = configurationMemory_io_out_bits_confneuralNetsbiasVecs_0_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVecs_0_1 = configurationMemory_io_out_bits_confneuralNetsbiasVecs_0_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVecs_0_2 = configurationMemory_io_out_bits_confneuralNetsbiasVecs_0_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVecs_0_3 = configurationMemory_io_out_bits_confneuralNetsbiasVecs_0_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVecs_0_4 = configurationMemory_io_out_bits_confneuralNetsbiasVecs_0_4; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVecs_0_5 = configurationMemory_io_out_bits_confneuralNetsbiasVecs_0_5; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVecs_0_6 = configurationMemory_io_out_bits_confneuralNetsbiasVecs_0_6; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVecs_0_7 = configurationMemory_io_out_bits_confneuralNetsbiasVecs_0_7; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVecs_0_8 = configurationMemory_io_out_bits_confneuralNetsbiasVecs_0_8; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVecs_0_9 = configurationMemory_io_out_bits_confneuralNetsbiasVecs_0_9; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVecs_1_0 = configurationMemory_io_out_bits_confneuralNetsbiasVecs_1_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVecs_1_1 = configurationMemory_io_out_bits_confneuralNetsbiasVecs_1_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVecs_1_2 = configurationMemory_io_out_bits_confneuralNetsbiasVecs_1_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVecs_1_3 = configurationMemory_io_out_bits_confneuralNetsbiasVecs_1_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVecs_1_4 = configurationMemory_io_out_bits_confneuralNetsbiasVecs_1_4; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVecs_1_5 = configurationMemory_io_out_bits_confneuralNetsbiasVecs_1_5; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVecs_1_6 = configurationMemory_io_out_bits_confneuralNetsbiasVecs_1_6; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVecs_1_7 = configurationMemory_io_out_bits_confneuralNetsbiasVecs_1_7; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVecs_1_8 = configurationMemory_io_out_bits_confneuralNetsbiasVecs_1_8; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVecs_1_9 = configurationMemory_io_out_bits_confneuralNetsbiasVecs_1_9; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVecs_2_0 = configurationMemory_io_out_bits_confneuralNetsbiasVecs_2_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVecs_2_1 = configurationMemory_io_out_bits_confneuralNetsbiasVecs_2_1; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVecs_2_2 = configurationMemory_io_out_bits_confneuralNetsbiasVecs_2_2; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVecs_2_3 = configurationMemory_io_out_bits_confneuralNetsbiasVecs_2_3; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVecs_2_4 = configurationMemory_io_out_bits_confneuralNetsbiasVecs_2_4; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVecs_2_5 = configurationMemory_io_out_bits_confneuralNetsbiasVecs_2_5; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVecs_2_6 = configurationMemory_io_out_bits_confneuralNetsbiasVecs_2_6; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVecs_2_7 = configurationMemory_io_out_bits_confneuralNetsbiasVecs_2_7; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVecs_2_8 = configurationMemory_io_out_bits_confneuralNetsbiasVecs_2_8; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsbiasVecs_2_9 = configurationMemory_io_out_bits_confneuralNetsbiasVecs_2_9; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confneuralNetsoutputBias_0 = configurationMemory_io_out_bits_confneuralNetsoutputBias_0; // @[Wellness.scala 420:24]
  assign wellness_io_inConf_bits_confInputMuxSel = configurationMemory_io_out_bits_confInputMuxSel; // @[Wellness.scala 420:24]
  assign configurationMemory_clock = clock;
  assign configurationMemory_reset = reset;
  assign configurationMemory_io_in_valid = converter_2_auto_out_valid; // @[Wellness.scala 416:37]
  assign configurationMemory_io_in_bits_wrdata = $signed(_T_7); // @[Wellness.scala 418:43]
  assign configurationMemory_io_in_bits_wraddr = inConf_bits_data[34:32]; // @[Wellness.scala 419:43]
endmodule
